-- floating_point.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity floating_point is
	port (
		clk_clk       : in  std_logic                     := '0';             --   clk.clk
		reset_reset_n : in  std_logic                     := '0';             -- reset.reset_n
		s1_dataa      : in  std_logic_vector(31 downto 0) := (others => '0'); --    s1.dataa
		s1_datab      : in  std_logic_vector(31 downto 0) := (others => '0'); --      .datab
		s1_n          : in  std_logic_vector(3 downto 0)  := (others => '0'); --      .n
		s1_result     : out std_logic_vector(31 downto 0);                    --      .result
		s2_clk        : in  std_logic                     := '0';             --    s2.clk
		s2_clk_en     : in  std_logic                     := '0';             --      .clk_en
		s2_dataa      : in  std_logic_vector(31 downto 0) := (others => '0'); --      .dataa
		s2_datab      : in  std_logic_vector(31 downto 0) := (others => '0'); --      .datab
		s2_n          : in  std_logic_vector(2 downto 0)  := (others => '0'); --      .n
		s2_reset      : in  std_logic                     := '0';             --      .reset
		s2_reset_req  : in  std_logic                     := '0';             --      .reset_req
		s2_start      : in  std_logic                     := '0';             --      .start
		s2_done       : out std_logic;                                        --      .done
		s2_result     : out std_logic_vector(31 downto 0)                     --      .result
	);
end entity floating_point;

architecture rtl of floating_point is
	component floating_point_nios_custom_instr_floating_point_2_0 is
		generic (
			sqrtf_enabled : integer := 1
		);
		port (
			s1_dataa     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			s1_datab     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			s1_n         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- n
			s1_result    : out std_logic_vector(31 downto 0);                    -- result
			s2_clk       : in  std_logic                     := 'X';             -- clk
			s2_clk_en    : in  std_logic                     := 'X';             -- clk_en
			s2_dataa     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			s2_datab     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			s2_n         : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- n
			s2_reset     : in  std_logic                     := 'X';             -- reset
			s2_reset_req : in  std_logic                     := 'X';             -- reset_req
			s2_start     : in  std_logic                     := 'X';             -- start
			s2_done      : out std_logic;                                        -- done
			s2_result    : out std_logic_vector(31 downto 0)                     -- result
		);
	end component floating_point_nios_custom_instr_floating_point_2_0;

begin

	nios_custom_instr_floating_point_2_0 : component floating_point_nios_custom_instr_floating_point_2_0
		generic map (
			sqrtf_enabled => 1
		)
		port map (
			s1_dataa     => s1_dataa,     -- s1.dataa
			s1_datab     => s1_datab,     --   .datab
			s1_n         => s1_n,         --   .n
			s1_result    => s1_result,    --   .result
			s2_clk       => s2_clk,       -- s2.clk
			s2_clk_en    => s2_clk_en,    --   .clk_en
			s2_dataa     => s2_dataa,     --   .dataa
			s2_datab     => s2_datab,     --   .datab
			s2_n         => s2_n,         --   .n
			s2_reset     => s2_reset,     --   .reset
			s2_reset_req => s2_reset_req, --   .reset_req
			s2_start     => s2_start,     --   .start
			s2_done      => s2_done,      --   .done
			s2_result    => s2_result     --   .result
		);

end architecture rtl; -- of floating_point
