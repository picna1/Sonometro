-- megafunction wizard: %ALTFP_LOG%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTFP_LOG 

-- ============================================================
-- File Name: prueba1.vhd
-- Megafunction Name(s):
-- 			ALTFP_LOG
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 15.1.0 Build 185 10/21/2015 SJ Lite Edition
-- ************************************************************


--Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, the Altera Quartus Prime License Agreement,
--the Altera MegaCore Function License Agreement, or other 
--applicable license agreement, including, without limitation, 
--that your use is for the sole purpose of programming logic 
--devices manufactured by Altera and sold by Altera or its 
--authorized distributors.  Please refer to the applicable 
--agreement for further details.


--altfp_log CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" PIPELINE=21 WIDTH_EXP=8 WIDTH_MAN=23 clock data result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" PIPELINE=1 SHIFTDIR="LEFT" WIDTH=32 WIDTHDIST=5 aclr clk_en clock data distance result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_mgl 2015:10:21:18:12:49:SJ  VERSION_END

--synthesis_resources = reg 33 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altbarrel_shift_05e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END prueba1_altbarrel_shift_05e;

 ARCHITECTURE RTL OF prueba1_altbarrel_shift_05e IS

	 SIGNAL	 dir_pipe	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper1d	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range264w276w277w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range264w272w273w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range285w297w298w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range285w293w294w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range307w319w320w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range307w315w316w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range329w341w342w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range329w337w338w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range351w363w364w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range351w359w360w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range264w268w269w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range285w289w290w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range307w311w312w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range329w333w334w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range351w355w356w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range264w276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range264w272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range285w297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range285w293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range307w319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range307w315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range329w341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range329w337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range351w363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range351w359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_dir_w_range261w275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_dir_w_range283w296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_dir_w_range304w318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_dir_w_range326w340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_dir_w_range348w362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range264w268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range285w289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range307w311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range329w333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_sel_w_range351w355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range264w276w277w278w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range285w297w298w299w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range307w319w320w321w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range329w341w342w343w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range351w363w364w365w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w279w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w300w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w322w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w344w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w366w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (191 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (159 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w271w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w274w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w292w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w295w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w314w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w317w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w336w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w339w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w358w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w361w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_dir_w_range261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_dir_w_range283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_dir_w_range304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_dir_w_range326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_dir_w_range348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sbit_w_range324w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sbit_w_range346w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sbit_w_range259w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sbit_w_range282w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sbit_w_range302w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sel_w_range264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sel_w_range285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sel_w_range307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sel_w_range329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_sel_w_range351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_w_smux_w_range367w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range264w276w277w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range264w276w(0) AND wire_Lshiftsmall_w274w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range264w272w273w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range264w272w(0) AND wire_Lshiftsmall_w271w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range285w297w298w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range285w297w(0) AND wire_Lshiftsmall_w295w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range285w293w294w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range285w293w(0) AND wire_Lshiftsmall_w292w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range307w319w320w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range307w319w(0) AND wire_Lshiftsmall_w317w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range307w315w316w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range307w315w(0) AND wire_Lshiftsmall_w314w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range329w341w342w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range329w341w(0) AND wire_Lshiftsmall_w339w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range329w337w338w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range329w337w(0) AND wire_Lshiftsmall_w336w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range351w363w364w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range351w363w(0) AND wire_Lshiftsmall_w361w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range351w359w360w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range351w359w(0) AND wire_Lshiftsmall_w358w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range264w268w269w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range264w268w(0) AND wire_Lshiftsmall_w_sbit_w_range259w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range285w289w290w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range285w289w(0) AND wire_Lshiftsmall_w_sbit_w_range282w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range307w311w312w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range307w311w(0) AND wire_Lshiftsmall_w_sbit_w_range302w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range329w333w334w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range329w333w(0) AND wire_Lshiftsmall_w_sbit_w_range324w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range351w355w356w(i) <= wire_Lshiftsmall_w_lg_w_sel_w_range351w355w(0) AND wire_Lshiftsmall_w_sbit_w_range346w(i);
	END GENERATE loop14;
	wire_Lshiftsmall_w_lg_w_sel_w_range264w276w(0) <= wire_Lshiftsmall_w_sel_w_range264w(0) AND wire_Lshiftsmall_w_lg_w_dir_w_range261w275w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range264w272w(0) <= wire_Lshiftsmall_w_sel_w_range264w(0) AND wire_Lshiftsmall_w_dir_w_range261w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range285w297w(0) <= wire_Lshiftsmall_w_sel_w_range285w(0) AND wire_Lshiftsmall_w_lg_w_dir_w_range283w296w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range285w293w(0) <= wire_Lshiftsmall_w_sel_w_range285w(0) AND wire_Lshiftsmall_w_dir_w_range283w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range307w319w(0) <= wire_Lshiftsmall_w_sel_w_range307w(0) AND wire_Lshiftsmall_w_lg_w_dir_w_range304w318w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range307w315w(0) <= wire_Lshiftsmall_w_sel_w_range307w(0) AND wire_Lshiftsmall_w_dir_w_range304w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range329w341w(0) <= wire_Lshiftsmall_w_sel_w_range329w(0) AND wire_Lshiftsmall_w_lg_w_dir_w_range326w340w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range329w337w(0) <= wire_Lshiftsmall_w_sel_w_range329w(0) AND wire_Lshiftsmall_w_dir_w_range326w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range351w363w(0) <= wire_Lshiftsmall_w_sel_w_range351w(0) AND wire_Lshiftsmall_w_lg_w_dir_w_range348w362w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range351w359w(0) <= wire_Lshiftsmall_w_sel_w_range351w(0) AND wire_Lshiftsmall_w_dir_w_range348w(0);
	wire_Lshiftsmall_w_lg_w_dir_w_range261w275w(0) <= NOT wire_Lshiftsmall_w_dir_w_range261w(0);
	wire_Lshiftsmall_w_lg_w_dir_w_range283w296w(0) <= NOT wire_Lshiftsmall_w_dir_w_range283w(0);
	wire_Lshiftsmall_w_lg_w_dir_w_range304w318w(0) <= NOT wire_Lshiftsmall_w_dir_w_range304w(0);
	wire_Lshiftsmall_w_lg_w_dir_w_range326w340w(0) <= NOT wire_Lshiftsmall_w_dir_w_range326w(0);
	wire_Lshiftsmall_w_lg_w_dir_w_range348w362w(0) <= NOT wire_Lshiftsmall_w_dir_w_range348w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range264w268w(0) <= NOT wire_Lshiftsmall_w_sel_w_range264w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range285w289w(0) <= NOT wire_Lshiftsmall_w_sel_w_range285w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range307w311w(0) <= NOT wire_Lshiftsmall_w_sel_w_range307w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range329w333w(0) <= NOT wire_Lshiftsmall_w_sel_w_range329w(0);
	wire_Lshiftsmall_w_lg_w_sel_w_range351w355w(0) <= NOT wire_Lshiftsmall_w_sel_w_range351w(0);
	loop15 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range264w276w277w278w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range264w276w277w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range264w272w273w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range285w297w298w299w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range285w297w298w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range285w293w294w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range307w319w320w321w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range307w319w320w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range307w315w316w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range329w341w342w343w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range329w341w342w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range329w337w338w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range351w363w364w365w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range351w363w364w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range351w359w360w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w279w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range264w276w277w278w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range264w268w269w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w300w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range285w297w298w299w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range285w289w290w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w322w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range307w319w320w321w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range307w311w312w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w344w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range329w341w342w343w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range329w333w334w(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 31 GENERATE 
		wire_Lshiftsmall_w366w(i) <= wire_Lshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range351w363w364w365w(i) OR wire_Lshiftsmall_w_lg_w_lg_w_sel_w_range351w355w356w(i);
	END GENERATE loop24;
	dir_w <= ( dir_pipe(0) & dir_w(3 DOWNTO 0) & direction_w);
	direction_w <= '0';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(191 DOWNTO 160);
	sbit_w <= ( sbit_piper1d & smux_w(127 DOWNTO 0) & data);
	sel_w <= ( distance(4 DOWNTO 0));
	smux_w <= ( wire_Lshiftsmall_w366w & wire_Lshiftsmall_w344w & wire_Lshiftsmall_w322w & wire_Lshiftsmall_w300w & wire_Lshiftsmall_w279w);
	wire_Lshiftsmall_w271w <= ( pad_w(0) & sbit_w(31 DOWNTO 1));
	wire_Lshiftsmall_w274w <= ( sbit_w(30 DOWNTO 0) & pad_w(0));
	wire_Lshiftsmall_w292w <= ( pad_w(1 DOWNTO 0) & sbit_w(63 DOWNTO 34));
	wire_Lshiftsmall_w295w <= ( sbit_w(61 DOWNTO 32) & pad_w(1 DOWNTO 0));
	wire_Lshiftsmall_w314w <= ( pad_w(3 DOWNTO 0) & sbit_w(95 DOWNTO 68));
	wire_Lshiftsmall_w317w <= ( sbit_w(91 DOWNTO 64) & pad_w(3 DOWNTO 0));
	wire_Lshiftsmall_w336w <= ( pad_w(7 DOWNTO 0) & sbit_w(127 DOWNTO 104));
	wire_Lshiftsmall_w339w <= ( sbit_w(119 DOWNTO 96) & pad_w(7 DOWNTO 0));
	wire_Lshiftsmall_w358w <= ( pad_w(15 DOWNTO 0) & sbit_w(159 DOWNTO 144));
	wire_Lshiftsmall_w361w <= ( sbit_w(143 DOWNTO 128) & pad_w(15 DOWNTO 0));
	wire_Lshiftsmall_w_dir_w_range261w(0) <= dir_w(0);
	wire_Lshiftsmall_w_dir_w_range283w(0) <= dir_w(1);
	wire_Lshiftsmall_w_dir_w_range304w(0) <= dir_w(2);
	wire_Lshiftsmall_w_dir_w_range326w(0) <= dir_w(3);
	wire_Lshiftsmall_w_dir_w_range348w(0) <= dir_w(4);
	wire_Lshiftsmall_w_sbit_w_range324w <= sbit_w(127 DOWNTO 96);
	wire_Lshiftsmall_w_sbit_w_range346w <= sbit_w(159 DOWNTO 128);
	wire_Lshiftsmall_w_sbit_w_range259w <= sbit_w(31 DOWNTO 0);
	wire_Lshiftsmall_w_sbit_w_range282w <= sbit_w(63 DOWNTO 32);
	wire_Lshiftsmall_w_sbit_w_range302w <= sbit_w(95 DOWNTO 64);
	wire_Lshiftsmall_w_sel_w_range264w(0) <= sel_w(0);
	wire_Lshiftsmall_w_sel_w_range285w(0) <= sel_w(1);
	wire_Lshiftsmall_w_sel_w_range307w(0) <= sel_w(2);
	wire_Lshiftsmall_w_sel_w_range329w(0) <= sel_w(3);
	wire_Lshiftsmall_w_sel_w_range351w(0) <= sel_w(4);
	wire_Lshiftsmall_w_smux_w_range367w <= smux_w(159 DOWNTO 128);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dir_pipe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dir_pipe(0) <= ( dir_w(4));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper1d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper1d <= wire_Lshiftsmall_w_smux_w_range367w;
			END IF;
		END IF;
	END PROCESS;

 END RTL; --prueba1_altbarrel_shift_05e


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" SHIFTDIR="LEFT" WIDTH=64 WIDTHDIST=6 data distance result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_mgl 2015:10:21:18:12:49:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altbarrel_shift_8ib IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (5 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (63 DOWNTO 0)
	 ); 
 END prueba1_altbarrel_shift_8ib;

 ARCHITECTURE RTL OF prueba1_altbarrel_shift_8ib IS

	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range378w390w391w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range378w386w387w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range399w411w412w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range399w407w408w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range421w433w434w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range421w429w430w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range443w455w456w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range443w451w452w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range465w477w478w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range465w473w474w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range487w499w500w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range487w495w496w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range378w382w383w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range399w403w404w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range421w425w426w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range443w447w448w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range465w469w470w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range487w491w492w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range378w390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range378w386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range399w411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range399w407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range421w433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range421w429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range443w455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range443w451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range465w477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range465w473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range487w499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range487w495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_dir_w_range375w389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_dir_w_range397w410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_dir_w_range418w432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_dir_w_range440w454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_dir_w_range462w476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_dir_w_range484w498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range378w382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range399w403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range421w425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range443w447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range465w469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_sel_w_range487w491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range378w390w391w392w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range399w411w412w413w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range421w433w434w435w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range443w455w456w457w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range465w477w478w479w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range487w499w500w501w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w393w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w414w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w436w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w458w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w480w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w502w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (447 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (383 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w385w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w388w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w406w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w409w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w428w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w431w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w450w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w453w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w472w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w475w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w494w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w497w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_dir_w_range375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_dir_w_range397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_dir_w_range418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_dir_w_range440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_dir_w_range462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_dir_w_range484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sbit_w_range396w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sbit_w_range416w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sbit_w_range438w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sbit_w_range460w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sbit_w_range482w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sbit_w_range373w	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sel_w_range378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sel_w_range399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sel_w_range421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sel_w_range443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sel_w_range465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_w_sel_w_range487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	loop25 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range378w390w391w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range378w390w(0) AND wire_lzc_norm_L_w388w(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range378w386w387w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range378w386w(0) AND wire_lzc_norm_L_w385w(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range399w411w412w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range399w411w(0) AND wire_lzc_norm_L_w409w(i);
	END GENERATE loop27;
	loop28 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range399w407w408w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range399w407w(0) AND wire_lzc_norm_L_w406w(i);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range421w433w434w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range421w433w(0) AND wire_lzc_norm_L_w431w(i);
	END GENERATE loop29;
	loop30 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range421w429w430w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range421w429w(0) AND wire_lzc_norm_L_w428w(i);
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range443w455w456w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range443w455w(0) AND wire_lzc_norm_L_w453w(i);
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range443w451w452w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range443w451w(0) AND wire_lzc_norm_L_w450w(i);
	END GENERATE loop32;
	loop33 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range465w477w478w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range465w477w(0) AND wire_lzc_norm_L_w475w(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range465w473w474w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range465w473w(0) AND wire_lzc_norm_L_w472w(i);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range487w499w500w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range487w499w(0) AND wire_lzc_norm_L_w497w(i);
	END GENERATE loop35;
	loop36 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range487w495w496w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range487w495w(0) AND wire_lzc_norm_L_w494w(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range378w382w383w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range378w382w(0) AND wire_lzc_norm_L_w_sbit_w_range373w(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range399w403w404w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range399w403w(0) AND wire_lzc_norm_L_w_sbit_w_range396w(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range421w425w426w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range421w425w(0) AND wire_lzc_norm_L_w_sbit_w_range416w(i);
	END GENERATE loop39;
	loop40 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range443w447w448w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range443w447w(0) AND wire_lzc_norm_L_w_sbit_w_range438w(i);
	END GENERATE loop40;
	loop41 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range465w469w470w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range465w469w(0) AND wire_lzc_norm_L_w_sbit_w_range460w(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range487w491w492w(i) <= wire_lzc_norm_L_w_lg_w_sel_w_range487w491w(0) AND wire_lzc_norm_L_w_sbit_w_range482w(i);
	END GENERATE loop42;
	wire_lzc_norm_L_w_lg_w_sel_w_range378w390w(0) <= wire_lzc_norm_L_w_sel_w_range378w(0) AND wire_lzc_norm_L_w_lg_w_dir_w_range375w389w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range378w386w(0) <= wire_lzc_norm_L_w_sel_w_range378w(0) AND wire_lzc_norm_L_w_dir_w_range375w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range399w411w(0) <= wire_lzc_norm_L_w_sel_w_range399w(0) AND wire_lzc_norm_L_w_lg_w_dir_w_range397w410w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range399w407w(0) <= wire_lzc_norm_L_w_sel_w_range399w(0) AND wire_lzc_norm_L_w_dir_w_range397w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range421w433w(0) <= wire_lzc_norm_L_w_sel_w_range421w(0) AND wire_lzc_norm_L_w_lg_w_dir_w_range418w432w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range421w429w(0) <= wire_lzc_norm_L_w_sel_w_range421w(0) AND wire_lzc_norm_L_w_dir_w_range418w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range443w455w(0) <= wire_lzc_norm_L_w_sel_w_range443w(0) AND wire_lzc_norm_L_w_lg_w_dir_w_range440w454w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range443w451w(0) <= wire_lzc_norm_L_w_sel_w_range443w(0) AND wire_lzc_norm_L_w_dir_w_range440w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range465w477w(0) <= wire_lzc_norm_L_w_sel_w_range465w(0) AND wire_lzc_norm_L_w_lg_w_dir_w_range462w476w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range465w473w(0) <= wire_lzc_norm_L_w_sel_w_range465w(0) AND wire_lzc_norm_L_w_dir_w_range462w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range487w499w(0) <= wire_lzc_norm_L_w_sel_w_range487w(0) AND wire_lzc_norm_L_w_lg_w_dir_w_range484w498w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range487w495w(0) <= wire_lzc_norm_L_w_sel_w_range487w(0) AND wire_lzc_norm_L_w_dir_w_range484w(0);
	wire_lzc_norm_L_w_lg_w_dir_w_range375w389w(0) <= NOT wire_lzc_norm_L_w_dir_w_range375w(0);
	wire_lzc_norm_L_w_lg_w_dir_w_range397w410w(0) <= NOT wire_lzc_norm_L_w_dir_w_range397w(0);
	wire_lzc_norm_L_w_lg_w_dir_w_range418w432w(0) <= NOT wire_lzc_norm_L_w_dir_w_range418w(0);
	wire_lzc_norm_L_w_lg_w_dir_w_range440w454w(0) <= NOT wire_lzc_norm_L_w_dir_w_range440w(0);
	wire_lzc_norm_L_w_lg_w_dir_w_range462w476w(0) <= NOT wire_lzc_norm_L_w_dir_w_range462w(0);
	wire_lzc_norm_L_w_lg_w_dir_w_range484w498w(0) <= NOT wire_lzc_norm_L_w_dir_w_range484w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range378w382w(0) <= NOT wire_lzc_norm_L_w_sel_w_range378w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range399w403w(0) <= NOT wire_lzc_norm_L_w_sel_w_range399w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range421w425w(0) <= NOT wire_lzc_norm_L_w_sel_w_range421w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range443w447w(0) <= NOT wire_lzc_norm_L_w_sel_w_range443w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range465w469w(0) <= NOT wire_lzc_norm_L_w_sel_w_range465w(0);
	wire_lzc_norm_L_w_lg_w_sel_w_range487w491w(0) <= NOT wire_lzc_norm_L_w_sel_w_range487w(0);
	loop43 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range378w390w391w392w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range378w390w391w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range378w386w387w(i);
	END GENERATE loop43;
	loop44 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range399w411w412w413w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range399w411w412w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range399w407w408w(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range421w433w434w435w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range421w433w434w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range421w429w430w(i);
	END GENERATE loop45;
	loop46 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range443w455w456w457w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range443w455w456w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range443w451w452w(i);
	END GENERATE loop46;
	loop47 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range465w477w478w479w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range465w477w478w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range465w473w474w(i);
	END GENERATE loop47;
	loop48 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range487w499w500w501w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range487w499w500w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range487w495w496w(i);
	END GENERATE loop48;
	loop49 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w393w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range378w390w391w392w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range378w382w383w(i);
	END GENERATE loop49;
	loop50 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w414w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range399w411w412w413w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range399w403w404w(i);
	END GENERATE loop50;
	loop51 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w436w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range421w433w434w435w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range421w425w426w(i);
	END GENERATE loop51;
	loop52 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w458w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range443w455w456w457w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range443w447w448w(i);
	END GENERATE loop52;
	loop53 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w480w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range465w477w478w479w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range465w469w470w(i);
	END GENERATE loop53;
	loop54 : FOR i IN 0 TO 63 GENERATE 
		wire_lzc_norm_L_w502w(i) <= wire_lzc_norm_L_w_lg_w_lg_w_lg_w_sel_w_range487w499w500w501w(i) OR wire_lzc_norm_L_w_lg_w_lg_w_sel_w_range487w491w492w(i);
	END GENERATE loop54;
	dir_w <= ( dir_w(5 DOWNTO 0) & direction_w);
	direction_w <= '0';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(447 DOWNTO 384);
	sbit_w <= ( smux_w(383 DOWNTO 0) & data);
	sel_w <= ( distance(5 DOWNTO 0));
	smux_w <= ( wire_lzc_norm_L_w502w & wire_lzc_norm_L_w480w & wire_lzc_norm_L_w458w & wire_lzc_norm_L_w436w & wire_lzc_norm_L_w414w & wire_lzc_norm_L_w393w);
	wire_lzc_norm_L_w385w <= ( pad_w(0) & sbit_w(63 DOWNTO 1));
	wire_lzc_norm_L_w388w <= ( sbit_w(62 DOWNTO 0) & pad_w(0));
	wire_lzc_norm_L_w406w <= ( pad_w(1 DOWNTO 0) & sbit_w(127 DOWNTO 66));
	wire_lzc_norm_L_w409w <= ( sbit_w(125 DOWNTO 64) & pad_w(1 DOWNTO 0));
	wire_lzc_norm_L_w428w <= ( pad_w(3 DOWNTO 0) & sbit_w(191 DOWNTO 132));
	wire_lzc_norm_L_w431w <= ( sbit_w(187 DOWNTO 128) & pad_w(3 DOWNTO 0));
	wire_lzc_norm_L_w450w <= ( pad_w(7 DOWNTO 0) & sbit_w(255 DOWNTO 200));
	wire_lzc_norm_L_w453w <= ( sbit_w(247 DOWNTO 192) & pad_w(7 DOWNTO 0));
	wire_lzc_norm_L_w472w <= ( pad_w(15 DOWNTO 0) & sbit_w(319 DOWNTO 272));
	wire_lzc_norm_L_w475w <= ( sbit_w(303 DOWNTO 256) & pad_w(15 DOWNTO 0));
	wire_lzc_norm_L_w494w <= ( pad_w(31 DOWNTO 0) & sbit_w(383 DOWNTO 352));
	wire_lzc_norm_L_w497w <= ( sbit_w(351 DOWNTO 320) & pad_w(31 DOWNTO 0));
	wire_lzc_norm_L_w_dir_w_range375w(0) <= dir_w(0);
	wire_lzc_norm_L_w_dir_w_range397w(0) <= dir_w(1);
	wire_lzc_norm_L_w_dir_w_range418w(0) <= dir_w(2);
	wire_lzc_norm_L_w_dir_w_range440w(0) <= dir_w(3);
	wire_lzc_norm_L_w_dir_w_range462w(0) <= dir_w(4);
	wire_lzc_norm_L_w_dir_w_range484w(0) <= dir_w(5);
	wire_lzc_norm_L_w_sbit_w_range396w <= sbit_w(127 DOWNTO 64);
	wire_lzc_norm_L_w_sbit_w_range416w <= sbit_w(191 DOWNTO 128);
	wire_lzc_norm_L_w_sbit_w_range438w <= sbit_w(255 DOWNTO 192);
	wire_lzc_norm_L_w_sbit_w_range460w <= sbit_w(319 DOWNTO 256);
	wire_lzc_norm_L_w_sbit_w_range482w <= sbit_w(383 DOWNTO 320);
	wire_lzc_norm_L_w_sbit_w_range373w <= sbit_w(63 DOWNTO 0);
	wire_lzc_norm_L_w_sel_w_range378w(0) <= sel_w(0);
	wire_lzc_norm_L_w_sel_w_range399w(0) <= sel_w(1);
	wire_lzc_norm_L_w_sel_w_range421w(0) <= sel_w(2);
	wire_lzc_norm_L_w_sel_w_range443w(0) <= sel_w(3);
	wire_lzc_norm_L_w_sel_w_range465w(0) <= sel_w(4);
	wire_lzc_norm_L_w_sel_w_range487w(0) <= sel_w(5);

 END RTL; --prueba1_altbarrel_shift_8ib


--altbarrel_shift CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" PIPELINE=1 SHIFTDIR="RIGHT" WIDTH=32 WIDTHDIST=5 aclr clk_en clock data distance result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_mgl 2015:10:21:18:12:49:SJ  VERSION_END

--synthesis_resources = reg 33 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altbarrel_shift_j8e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 distance	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END prueba1_altbarrel_shift_j8e;

 ARCHITECTURE RTL OF prueba1_altbarrel_shift_j8e IS

	 SIGNAL	 dir_pipe	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sbit_piper1d	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range514w526w527w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range514w522w523w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range535w547w548w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range535w543w544w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range557w569w570w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range557w565w566w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range579w591w592w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range579w587w588w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range601w613w614w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range601w609w610w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range514w518w519w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range535w539w540w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range557w561w562w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range579w583w584w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range601w605w606w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range514w526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range514w522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range535w547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range535w543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range557w569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range557w565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range579w591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range579w587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range601w613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range601w609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_dir_w_range511w525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_dir_w_range533w546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_dir_w_range554w568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_dir_w_range576w590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_dir_w_range598w612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range514w518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range535w539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range557w561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range579w583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_sel_w_range601w605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range514w526w527w528w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range535w547w548w549w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range557w569w570w571w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range579w591w592w593w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range601w613w614w615w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w529w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w550w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w572w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w594w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w616w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  dir_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  direction_w :	STD_LOGIC;
	 SIGNAL  pad_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  sbit_w :	STD_LOGIC_VECTOR (191 DOWNTO 0);
	 SIGNAL  sel_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  smux_w :	STD_LOGIC_VECTOR (159 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w521w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w524w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w542w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w545w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w564w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w567w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w586w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w589w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w608w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w611w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_dir_w_range511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_dir_w_range533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_dir_w_range554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_dir_w_range576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_dir_w_range598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sbit_w_range574w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sbit_w_range596w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sbit_w_range509w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sbit_w_range532w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sbit_w_range552w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sel_w_range514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sel_w_range535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sel_w_range557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sel_w_range579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_sel_w_range601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_w_smux_w_range617w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop55 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range514w526w527w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range514w526w(0) AND wire_Rshiftsmall_w524w(i);
	END GENERATE loop55;
	loop56 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range514w522w523w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range514w522w(0) AND wire_Rshiftsmall_w521w(i);
	END GENERATE loop56;
	loop57 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range535w547w548w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range535w547w(0) AND wire_Rshiftsmall_w545w(i);
	END GENERATE loop57;
	loop58 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range535w543w544w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range535w543w(0) AND wire_Rshiftsmall_w542w(i);
	END GENERATE loop58;
	loop59 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range557w569w570w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range557w569w(0) AND wire_Rshiftsmall_w567w(i);
	END GENERATE loop59;
	loop60 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range557w565w566w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range557w565w(0) AND wire_Rshiftsmall_w564w(i);
	END GENERATE loop60;
	loop61 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range579w591w592w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range579w591w(0) AND wire_Rshiftsmall_w589w(i);
	END GENERATE loop61;
	loop62 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range579w587w588w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range579w587w(0) AND wire_Rshiftsmall_w586w(i);
	END GENERATE loop62;
	loop63 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range601w613w614w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range601w613w(0) AND wire_Rshiftsmall_w611w(i);
	END GENERATE loop63;
	loop64 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range601w609w610w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range601w609w(0) AND wire_Rshiftsmall_w608w(i);
	END GENERATE loop64;
	loop65 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range514w518w519w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range514w518w(0) AND wire_Rshiftsmall_w_sbit_w_range509w(i);
	END GENERATE loop65;
	loop66 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range535w539w540w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range535w539w(0) AND wire_Rshiftsmall_w_sbit_w_range532w(i);
	END GENERATE loop66;
	loop67 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range557w561w562w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range557w561w(0) AND wire_Rshiftsmall_w_sbit_w_range552w(i);
	END GENERATE loop67;
	loop68 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range579w583w584w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range579w583w(0) AND wire_Rshiftsmall_w_sbit_w_range574w(i);
	END GENERATE loop68;
	loop69 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range601w605w606w(i) <= wire_Rshiftsmall_w_lg_w_sel_w_range601w605w(0) AND wire_Rshiftsmall_w_sbit_w_range596w(i);
	END GENERATE loop69;
	wire_Rshiftsmall_w_lg_w_sel_w_range514w526w(0) <= wire_Rshiftsmall_w_sel_w_range514w(0) AND wire_Rshiftsmall_w_lg_w_dir_w_range511w525w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range514w522w(0) <= wire_Rshiftsmall_w_sel_w_range514w(0) AND wire_Rshiftsmall_w_dir_w_range511w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range535w547w(0) <= wire_Rshiftsmall_w_sel_w_range535w(0) AND wire_Rshiftsmall_w_lg_w_dir_w_range533w546w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range535w543w(0) <= wire_Rshiftsmall_w_sel_w_range535w(0) AND wire_Rshiftsmall_w_dir_w_range533w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range557w569w(0) <= wire_Rshiftsmall_w_sel_w_range557w(0) AND wire_Rshiftsmall_w_lg_w_dir_w_range554w568w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range557w565w(0) <= wire_Rshiftsmall_w_sel_w_range557w(0) AND wire_Rshiftsmall_w_dir_w_range554w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range579w591w(0) <= wire_Rshiftsmall_w_sel_w_range579w(0) AND wire_Rshiftsmall_w_lg_w_dir_w_range576w590w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range579w587w(0) <= wire_Rshiftsmall_w_sel_w_range579w(0) AND wire_Rshiftsmall_w_dir_w_range576w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range601w613w(0) <= wire_Rshiftsmall_w_sel_w_range601w(0) AND wire_Rshiftsmall_w_lg_w_dir_w_range598w612w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range601w609w(0) <= wire_Rshiftsmall_w_sel_w_range601w(0) AND wire_Rshiftsmall_w_dir_w_range598w(0);
	wire_Rshiftsmall_w_lg_w_dir_w_range511w525w(0) <= NOT wire_Rshiftsmall_w_dir_w_range511w(0);
	wire_Rshiftsmall_w_lg_w_dir_w_range533w546w(0) <= NOT wire_Rshiftsmall_w_dir_w_range533w(0);
	wire_Rshiftsmall_w_lg_w_dir_w_range554w568w(0) <= NOT wire_Rshiftsmall_w_dir_w_range554w(0);
	wire_Rshiftsmall_w_lg_w_dir_w_range576w590w(0) <= NOT wire_Rshiftsmall_w_dir_w_range576w(0);
	wire_Rshiftsmall_w_lg_w_dir_w_range598w612w(0) <= NOT wire_Rshiftsmall_w_dir_w_range598w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range514w518w(0) <= NOT wire_Rshiftsmall_w_sel_w_range514w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range535w539w(0) <= NOT wire_Rshiftsmall_w_sel_w_range535w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range557w561w(0) <= NOT wire_Rshiftsmall_w_sel_w_range557w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range579w583w(0) <= NOT wire_Rshiftsmall_w_sel_w_range579w(0);
	wire_Rshiftsmall_w_lg_w_sel_w_range601w605w(0) <= NOT wire_Rshiftsmall_w_sel_w_range601w(0);
	loop70 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range514w526w527w528w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range514w526w527w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range514w522w523w(i);
	END GENERATE loop70;
	loop71 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range535w547w548w549w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range535w547w548w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range535w543w544w(i);
	END GENERATE loop71;
	loop72 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range557w569w570w571w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range557w569w570w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range557w565w566w(i);
	END GENERATE loop72;
	loop73 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range579w591w592w593w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range579w591w592w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range579w587w588w(i);
	END GENERATE loop73;
	loop74 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range601w613w614w615w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range601w613w614w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range601w609w610w(i);
	END GENERATE loop74;
	loop75 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w529w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range514w526w527w528w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range514w518w519w(i);
	END GENERATE loop75;
	loop76 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w550w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range535w547w548w549w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range535w539w540w(i);
	END GENERATE loop76;
	loop77 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w572w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range557w569w570w571w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range557w561w562w(i);
	END GENERATE loop77;
	loop78 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w594w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range579w591w592w593w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range579w583w584w(i);
	END GENERATE loop78;
	loop79 : FOR i IN 0 TO 31 GENERATE 
		wire_Rshiftsmall_w616w(i) <= wire_Rshiftsmall_w_lg_w_lg_w_lg_w_sel_w_range601w613w614w615w(i) OR wire_Rshiftsmall_w_lg_w_lg_w_sel_w_range601w605w606w(i);
	END GENERATE loop79;
	dir_w <= ( dir_pipe(0) & dir_w(3 DOWNTO 0) & direction_w);
	direction_w <= '1';
	pad_w <= (OTHERS => '0');
	result <= sbit_w(191 DOWNTO 160);
	sbit_w <= ( sbit_piper1d & smux_w(127 DOWNTO 0) & data);
	sel_w <= ( distance(4 DOWNTO 0));
	smux_w <= ( wire_Rshiftsmall_w616w & wire_Rshiftsmall_w594w & wire_Rshiftsmall_w572w & wire_Rshiftsmall_w550w & wire_Rshiftsmall_w529w);
	wire_Rshiftsmall_w521w <= ( pad_w(0) & sbit_w(31 DOWNTO 1));
	wire_Rshiftsmall_w524w <= ( sbit_w(30 DOWNTO 0) & pad_w(0));
	wire_Rshiftsmall_w542w <= ( pad_w(1 DOWNTO 0) & sbit_w(63 DOWNTO 34));
	wire_Rshiftsmall_w545w <= ( sbit_w(61 DOWNTO 32) & pad_w(1 DOWNTO 0));
	wire_Rshiftsmall_w564w <= ( pad_w(3 DOWNTO 0) & sbit_w(95 DOWNTO 68));
	wire_Rshiftsmall_w567w <= ( sbit_w(91 DOWNTO 64) & pad_w(3 DOWNTO 0));
	wire_Rshiftsmall_w586w <= ( pad_w(7 DOWNTO 0) & sbit_w(127 DOWNTO 104));
	wire_Rshiftsmall_w589w <= ( sbit_w(119 DOWNTO 96) & pad_w(7 DOWNTO 0));
	wire_Rshiftsmall_w608w <= ( pad_w(15 DOWNTO 0) & sbit_w(159 DOWNTO 144));
	wire_Rshiftsmall_w611w <= ( sbit_w(143 DOWNTO 128) & pad_w(15 DOWNTO 0));
	wire_Rshiftsmall_w_dir_w_range511w(0) <= dir_w(0);
	wire_Rshiftsmall_w_dir_w_range533w(0) <= dir_w(1);
	wire_Rshiftsmall_w_dir_w_range554w(0) <= dir_w(2);
	wire_Rshiftsmall_w_dir_w_range576w(0) <= dir_w(3);
	wire_Rshiftsmall_w_dir_w_range598w(0) <= dir_w(4);
	wire_Rshiftsmall_w_sbit_w_range574w <= sbit_w(127 DOWNTO 96);
	wire_Rshiftsmall_w_sbit_w_range596w <= sbit_w(159 DOWNTO 128);
	wire_Rshiftsmall_w_sbit_w_range509w <= sbit_w(31 DOWNTO 0);
	wire_Rshiftsmall_w_sbit_w_range532w <= sbit_w(63 DOWNTO 32);
	wire_Rshiftsmall_w_sbit_w_range552w <= sbit_w(95 DOWNTO 64);
	wire_Rshiftsmall_w_sel_w_range514w(0) <= sel_w(0);
	wire_Rshiftsmall_w_sel_w_range535w(0) <= sel_w(1);
	wire_Rshiftsmall_w_sel_w_range557w(0) <= sel_w(2);
	wire_Rshiftsmall_w_sel_w_range579w(0) <= sel_w(3);
	wire_Rshiftsmall_w_sel_w_range601w(0) <= sel_w(4);
	wire_Rshiftsmall_w_smux_w_range617w <= smux_w(159 DOWNTO 128);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN dir_pipe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN dir_pipe(0) <= ( dir_w(4));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sbit_piper1d <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sbit_piper1d <= wire_Rshiftsmall_w_smux_w_range617w;
			END IF;
		END IF;
	END PROCESS;

 END RTL; --prueba1_altbarrel_shift_j8e


--altfp_log_and_or CBX_AUTO_BLACKBOX="ALL" LUT_INPUT_COUNT=4 OPERATION="AND" PIPELINE=3 WIDTH=8 aclr clken clock data result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

--synthesis_resources = reg 4 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_and_or_f9b IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC
	 ); 
 END prueba1_altfp_log_and_or_f9b;

 ARCHITECTURE RTL OF prueba1_altfp_log_and_or_f9b IS

	 SIGNAL	 connection_dffe0	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exp_nan_w_lg_w_operation_r1_w_range624w628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_lg_w_operation_r1_w_range627w631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_lg_w_operation_r1_w_range630w634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_lg_w_operation_r1_w_range636w639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_lg_w_operation_r1_w_range638w642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_lg_w_operation_r1_w_range641w645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_lg_w_operation_r2_w_range651w655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  connection_r0_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  connection_r1_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  connection_r2_w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  operation_r1_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  operation_r2_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_connection_r0_w_range626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_connection_r0_w_range629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_connection_r0_w_range632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_connection_r0_w_range637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_connection_r0_w_range640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_connection_r0_w_range643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_connection_r1_w_range653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_operation_r1_w_range624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_operation_r1_w_range627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_operation_r1_w_range630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_operation_r1_w_range636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_operation_r1_w_range638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_operation_r1_w_range641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_nan_w_operation_r2_w_range651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_exp_nan_w_lg_w_operation_r1_w_range624w628w(0) <= wire_exp_nan_w_operation_r1_w_range624w(0) AND wire_exp_nan_w_connection_r0_w_range626w(0);
	wire_exp_nan_w_lg_w_operation_r1_w_range627w631w(0) <= wire_exp_nan_w_operation_r1_w_range627w(0) AND wire_exp_nan_w_connection_r0_w_range629w(0);
	wire_exp_nan_w_lg_w_operation_r1_w_range630w634w(0) <= wire_exp_nan_w_operation_r1_w_range630w(0) AND wire_exp_nan_w_connection_r0_w_range632w(0);
	wire_exp_nan_w_lg_w_operation_r1_w_range636w639w(0) <= wire_exp_nan_w_operation_r1_w_range636w(0) AND wire_exp_nan_w_connection_r0_w_range637w(0);
	wire_exp_nan_w_lg_w_operation_r1_w_range638w642w(0) <= wire_exp_nan_w_operation_r1_w_range638w(0) AND wire_exp_nan_w_connection_r0_w_range640w(0);
	wire_exp_nan_w_lg_w_operation_r1_w_range641w645w(0) <= wire_exp_nan_w_operation_r1_w_range641w(0) AND wire_exp_nan_w_connection_r0_w_range643w(0);
	wire_exp_nan_w_lg_w_operation_r2_w_range651w655w(0) <= wire_exp_nan_w_operation_r2_w_range651w(0) AND wire_exp_nan_w_connection_r1_w_range653w(0);
	connection_r0_w <= data;
	connection_r1_w <= connection_dffe0;
	connection_r2_w <= connection_dffe1;
	operation_r1_w <= ( wire_exp_nan_w_lg_w_operation_r1_w_range641w645w & wire_exp_nan_w_lg_w_operation_r1_w_range638w642w & wire_exp_nan_w_lg_w_operation_r1_w_range636w639w & connection_r0_w(4) & wire_exp_nan_w_lg_w_operation_r1_w_range630w634w & wire_exp_nan_w_lg_w_operation_r1_w_range627w631w & wire_exp_nan_w_lg_w_operation_r1_w_range624w628w & connection_r0_w(0));
	operation_r2_w <= ( wire_exp_nan_w_lg_w_operation_r2_w_range651w655w & connection_r1_w(0));
	result <= connection_dffe2;
	wire_exp_nan_w_connection_r0_w_range626w(0) <= connection_r0_w(1);
	wire_exp_nan_w_connection_r0_w_range629w(0) <= connection_r0_w(2);
	wire_exp_nan_w_connection_r0_w_range632w(0) <= connection_r0_w(3);
	wire_exp_nan_w_connection_r0_w_range637w(0) <= connection_r0_w(5);
	wire_exp_nan_w_connection_r0_w_range640w(0) <= connection_r0_w(6);
	wire_exp_nan_w_connection_r0_w_range643w(0) <= connection_r0_w(7);
	wire_exp_nan_w_connection_r1_w_range653w(0) <= connection_r1_w(1);
	wire_exp_nan_w_operation_r1_w_range624w(0) <= operation_r1_w(0);
	wire_exp_nan_w_operation_r1_w_range627w(0) <= operation_r1_w(1);
	wire_exp_nan_w_operation_r1_w_range630w(0) <= operation_r1_w(2);
	wire_exp_nan_w_operation_r1_w_range636w(0) <= operation_r1_w(4);
	wire_exp_nan_w_operation_r1_w_range638w(0) <= operation_r1_w(5);
	wire_exp_nan_w_operation_r1_w_range641w(0) <= operation_r1_w(6);
	wire_exp_nan_w_operation_r2_w_range651w(0) <= operation_r2_w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe0 <= ( operation_r1_w(7) & operation_r1_w(3));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe1(0) <= ( operation_r2_w(1));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe2 <= connection_r2_w(0);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --prueba1_altfp_log_and_or_f9b


--altfp_log_and_or CBX_AUTO_BLACKBOX="ALL" LUT_INPUT_COUNT=4 OPERATION="OR" PIPELINE=3 WIDTH=8 aclr clken clock data result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

--synthesis_resources = reg 4 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_and_or_t6b IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC
	 ); 
 END prueba1_altfp_log_and_or_t6b;

 ARCHITECTURE RTL OF prueba1_altfp_log_and_or_t6b IS

	 SIGNAL	 connection_dffe0	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exp_zero_w_lg_w_operation_r1_w_range660w664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_lg_w_operation_r1_w_range663w667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_lg_w_operation_r1_w_range666w670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_lg_w_operation_r1_w_range672w675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_lg_w_operation_r1_w_range674w678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_lg_w_operation_r1_w_range677w681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_lg_w_operation_r2_w_range687w691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  connection_r0_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  connection_r1_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  connection_r2_w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  operation_r1_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  operation_r2_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_connection_r0_w_range662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_connection_r0_w_range665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_connection_r0_w_range668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_connection_r0_w_range673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_connection_r0_w_range676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_connection_r0_w_range679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_connection_r1_w_range689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_operation_r1_w_range660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_operation_r1_w_range663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_operation_r1_w_range666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_operation_r1_w_range672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_operation_r1_w_range674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_operation_r1_w_range677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_zero_w_operation_r2_w_range687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_exp_zero_w_lg_w_operation_r1_w_range660w664w(0) <= wire_exp_zero_w_operation_r1_w_range660w(0) OR wire_exp_zero_w_connection_r0_w_range662w(0);
	wire_exp_zero_w_lg_w_operation_r1_w_range663w667w(0) <= wire_exp_zero_w_operation_r1_w_range663w(0) OR wire_exp_zero_w_connection_r0_w_range665w(0);
	wire_exp_zero_w_lg_w_operation_r1_w_range666w670w(0) <= wire_exp_zero_w_operation_r1_w_range666w(0) OR wire_exp_zero_w_connection_r0_w_range668w(0);
	wire_exp_zero_w_lg_w_operation_r1_w_range672w675w(0) <= wire_exp_zero_w_operation_r1_w_range672w(0) OR wire_exp_zero_w_connection_r0_w_range673w(0);
	wire_exp_zero_w_lg_w_operation_r1_w_range674w678w(0) <= wire_exp_zero_w_operation_r1_w_range674w(0) OR wire_exp_zero_w_connection_r0_w_range676w(0);
	wire_exp_zero_w_lg_w_operation_r1_w_range677w681w(0) <= wire_exp_zero_w_operation_r1_w_range677w(0) OR wire_exp_zero_w_connection_r0_w_range679w(0);
	wire_exp_zero_w_lg_w_operation_r2_w_range687w691w(0) <= wire_exp_zero_w_operation_r2_w_range687w(0) OR wire_exp_zero_w_connection_r1_w_range689w(0);
	connection_r0_w <= data;
	connection_r1_w <= connection_dffe0;
	connection_r2_w <= connection_dffe1;
	operation_r1_w <= ( wire_exp_zero_w_lg_w_operation_r1_w_range677w681w & wire_exp_zero_w_lg_w_operation_r1_w_range674w678w & wire_exp_zero_w_lg_w_operation_r1_w_range672w675w & connection_r0_w(4) & wire_exp_zero_w_lg_w_operation_r1_w_range666w670w & wire_exp_zero_w_lg_w_operation_r1_w_range663w667w & wire_exp_zero_w_lg_w_operation_r1_w_range660w664w & connection_r0_w(0));
	operation_r2_w <= ( wire_exp_zero_w_lg_w_operation_r2_w_range687w691w & connection_r1_w(0));
	result <= connection_dffe2;
	wire_exp_zero_w_connection_r0_w_range662w(0) <= connection_r0_w(1);
	wire_exp_zero_w_connection_r0_w_range665w(0) <= connection_r0_w(2);
	wire_exp_zero_w_connection_r0_w_range668w(0) <= connection_r0_w(3);
	wire_exp_zero_w_connection_r0_w_range673w(0) <= connection_r0_w(5);
	wire_exp_zero_w_connection_r0_w_range676w(0) <= connection_r0_w(6);
	wire_exp_zero_w_connection_r0_w_range679w(0) <= connection_r0_w(7);
	wire_exp_zero_w_connection_r1_w_range689w(0) <= connection_r1_w(1);
	wire_exp_zero_w_operation_r1_w_range660w(0) <= operation_r1_w(0);
	wire_exp_zero_w_operation_r1_w_range663w(0) <= operation_r1_w(1);
	wire_exp_zero_w_operation_r1_w_range666w(0) <= operation_r1_w(2);
	wire_exp_zero_w_operation_r1_w_range672w(0) <= operation_r1_w(4);
	wire_exp_zero_w_operation_r1_w_range674w(0) <= operation_r1_w(5);
	wire_exp_zero_w_operation_r1_w_range677w(0) <= operation_r1_w(6);
	wire_exp_zero_w_operation_r2_w_range687w(0) <= operation_r2_w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe0 <= ( operation_r1_w(7) & operation_r1_w(3));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe1(0) <= ( operation_r2_w(1));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe2 <= connection_r2_w(0);
			END IF;
		END IF;
	END PROCESS;

 END RTL; --prueba1_altfp_log_and_or_t6b


--altfp_log_and_or CBX_AUTO_BLACKBOX="ALL" LUT_INPUT_COUNT=4 OPERATION="OR" PIPELINE=3 WIDTH=23 aclr clken clock data result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

--synthesis_resources = reg 9 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_and_or_a8b IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (22 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC
	 ); 
 END prueba1_altfp_log_and_or_a8b;

 ARCHITECTURE RTL OF prueba1_altfp_log_and_or_a8b IS

	 SIGNAL	 connection_dffe0	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe1	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 connection_dffe2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range696w700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range724w728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range730w733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range732w736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range735w739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range741w744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range743w747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range746w750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range699w703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range752w755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range754w758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range702w706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range708w711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range710w714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range713w717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range719w722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r1_w_range721w725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r2_w_range768w772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r2_w_range771w775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r2_w_range774w778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r2_w_range780w783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_lg_w_operation_r3_w_range788w792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  connection_r0_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  connection_r1_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  connection_r2_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  connection_r3_w :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  operation_r1_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  operation_r2_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  operation_r3_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r0_w_range720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r1_w_range770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r1_w_range773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r1_w_range776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r1_w_range781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_connection_r2_w_range790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r1_w_range721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r2_w_range768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r2_w_range771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r2_w_range774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r2_w_range780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_inf_w_operation_r3_w_range788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
 BEGIN

	wire_man_inf_w_lg_w_operation_r1_w_range696w700w(0) <= wire_man_inf_w_operation_r1_w_range696w(0) OR wire_man_inf_w_connection_r0_w_range698w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range724w728w(0) <= wire_man_inf_w_operation_r1_w_range724w(0) OR wire_man_inf_w_connection_r0_w_range726w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range730w733w(0) <= wire_man_inf_w_operation_r1_w_range730w(0) OR wire_man_inf_w_connection_r0_w_range731w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range732w736w(0) <= wire_man_inf_w_operation_r1_w_range732w(0) OR wire_man_inf_w_connection_r0_w_range734w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range735w739w(0) <= wire_man_inf_w_operation_r1_w_range735w(0) OR wire_man_inf_w_connection_r0_w_range737w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range741w744w(0) <= wire_man_inf_w_operation_r1_w_range741w(0) OR wire_man_inf_w_connection_r0_w_range742w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range743w747w(0) <= wire_man_inf_w_operation_r1_w_range743w(0) OR wire_man_inf_w_connection_r0_w_range745w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range746w750w(0) <= wire_man_inf_w_operation_r1_w_range746w(0) OR wire_man_inf_w_connection_r0_w_range748w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range699w703w(0) <= wire_man_inf_w_operation_r1_w_range699w(0) OR wire_man_inf_w_connection_r0_w_range701w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range752w755w(0) <= wire_man_inf_w_operation_r1_w_range752w(0) OR wire_man_inf_w_connection_r0_w_range753w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range754w758w(0) <= wire_man_inf_w_operation_r1_w_range754w(0) OR wire_man_inf_w_connection_r0_w_range756w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range702w706w(0) <= wire_man_inf_w_operation_r1_w_range702w(0) OR wire_man_inf_w_connection_r0_w_range704w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range708w711w(0) <= wire_man_inf_w_operation_r1_w_range708w(0) OR wire_man_inf_w_connection_r0_w_range709w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range710w714w(0) <= wire_man_inf_w_operation_r1_w_range710w(0) OR wire_man_inf_w_connection_r0_w_range712w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range713w717w(0) <= wire_man_inf_w_operation_r1_w_range713w(0) OR wire_man_inf_w_connection_r0_w_range715w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range719w722w(0) <= wire_man_inf_w_operation_r1_w_range719w(0) OR wire_man_inf_w_connection_r0_w_range720w(0);
	wire_man_inf_w_lg_w_operation_r1_w_range721w725w(0) <= wire_man_inf_w_operation_r1_w_range721w(0) OR wire_man_inf_w_connection_r0_w_range723w(0);
	wire_man_inf_w_lg_w_operation_r2_w_range768w772w(0) <= wire_man_inf_w_operation_r2_w_range768w(0) OR wire_man_inf_w_connection_r1_w_range770w(0);
	wire_man_inf_w_lg_w_operation_r2_w_range771w775w(0) <= wire_man_inf_w_operation_r2_w_range771w(0) OR wire_man_inf_w_connection_r1_w_range773w(0);
	wire_man_inf_w_lg_w_operation_r2_w_range774w778w(0) <= wire_man_inf_w_operation_r2_w_range774w(0) OR wire_man_inf_w_connection_r1_w_range776w(0);
	wire_man_inf_w_lg_w_operation_r2_w_range780w783w(0) <= wire_man_inf_w_operation_r2_w_range780w(0) OR wire_man_inf_w_connection_r1_w_range781w(0);
	wire_man_inf_w_lg_w_operation_r3_w_range788w792w(0) <= wire_man_inf_w_operation_r3_w_range788w(0) OR wire_man_inf_w_connection_r2_w_range790w(0);
	connection_r0_w <= data;
	connection_r1_w <= connection_dffe0;
	connection_r2_w <= connection_dffe1;
	connection_r3_w <= connection_dffe2;
	operation_r1_w <= ( wire_man_inf_w_lg_w_operation_r1_w_range754w758w & wire_man_inf_w_lg_w_operation_r1_w_range752w755w & connection_r0_w(20) & wire_man_inf_w_lg_w_operation_r1_w_range746w750w & wire_man_inf_w_lg_w_operation_r1_w_range743w747w & wire_man_inf_w_lg_w_operation_r1_w_range741w744w & connection_r0_w(16) & wire_man_inf_w_lg_w_operation_r1_w_range735w739w & wire_man_inf_w_lg_w_operation_r1_w_range732w736w & wire_man_inf_w_lg_w_operation_r1_w_range730w733w & connection_r0_w(12) & wire_man_inf_w_lg_w_operation_r1_w_range724w728w & wire_man_inf_w_lg_w_operation_r1_w_range721w725w & wire_man_inf_w_lg_w_operation_r1_w_range719w722w & connection_r0_w(8) & wire_man_inf_w_lg_w_operation_r1_w_range713w717w & wire_man_inf_w_lg_w_operation_r1_w_range710w714w & wire_man_inf_w_lg_w_operation_r1_w_range708w711w & connection_r0_w(4) & wire_man_inf_w_lg_w_operation_r1_w_range702w706w & wire_man_inf_w_lg_w_operation_r1_w_range699w703w & wire_man_inf_w_lg_w_operation_r1_w_range696w700w & connection_r0_w(0));
	operation_r2_w <= ( wire_man_inf_w_lg_w_operation_r2_w_range780w783w & connection_r1_w(4) & wire_man_inf_w_lg_w_operation_r2_w_range774w778w & wire_man_inf_w_lg_w_operation_r2_w_range771w775w & wire_man_inf_w_lg_w_operation_r2_w_range768w772w & connection_r1_w(0));
	operation_r3_w <= ( wire_man_inf_w_lg_w_operation_r3_w_range788w792w & connection_r2_w(0));
	result <= connection_r3_w(0);
	wire_man_inf_w_connection_r0_w_range723w(0) <= connection_r0_w(10);
	wire_man_inf_w_connection_r0_w_range726w(0) <= connection_r0_w(11);
	wire_man_inf_w_connection_r0_w_range731w(0) <= connection_r0_w(13);
	wire_man_inf_w_connection_r0_w_range734w(0) <= connection_r0_w(14);
	wire_man_inf_w_connection_r0_w_range737w(0) <= connection_r0_w(15);
	wire_man_inf_w_connection_r0_w_range742w(0) <= connection_r0_w(17);
	wire_man_inf_w_connection_r0_w_range745w(0) <= connection_r0_w(18);
	wire_man_inf_w_connection_r0_w_range748w(0) <= connection_r0_w(19);
	wire_man_inf_w_connection_r0_w_range698w(0) <= connection_r0_w(1);
	wire_man_inf_w_connection_r0_w_range753w(0) <= connection_r0_w(21);
	wire_man_inf_w_connection_r0_w_range756w(0) <= connection_r0_w(22);
	wire_man_inf_w_connection_r0_w_range701w(0) <= connection_r0_w(2);
	wire_man_inf_w_connection_r0_w_range704w(0) <= connection_r0_w(3);
	wire_man_inf_w_connection_r0_w_range709w(0) <= connection_r0_w(5);
	wire_man_inf_w_connection_r0_w_range712w(0) <= connection_r0_w(6);
	wire_man_inf_w_connection_r0_w_range715w(0) <= connection_r0_w(7);
	wire_man_inf_w_connection_r0_w_range720w(0) <= connection_r0_w(9);
	wire_man_inf_w_connection_r1_w_range770w(0) <= connection_r1_w(1);
	wire_man_inf_w_connection_r1_w_range773w(0) <= connection_r1_w(2);
	wire_man_inf_w_connection_r1_w_range776w(0) <= connection_r1_w(3);
	wire_man_inf_w_connection_r1_w_range781w(0) <= connection_r1_w(5);
	wire_man_inf_w_connection_r2_w_range790w(0) <= connection_r2_w(1);
	wire_man_inf_w_operation_r1_w_range696w(0) <= operation_r1_w(0);
	wire_man_inf_w_operation_r1_w_range724w(0) <= operation_r1_w(10);
	wire_man_inf_w_operation_r1_w_range730w(0) <= operation_r1_w(12);
	wire_man_inf_w_operation_r1_w_range732w(0) <= operation_r1_w(13);
	wire_man_inf_w_operation_r1_w_range735w(0) <= operation_r1_w(14);
	wire_man_inf_w_operation_r1_w_range741w(0) <= operation_r1_w(16);
	wire_man_inf_w_operation_r1_w_range743w(0) <= operation_r1_w(17);
	wire_man_inf_w_operation_r1_w_range746w(0) <= operation_r1_w(18);
	wire_man_inf_w_operation_r1_w_range699w(0) <= operation_r1_w(1);
	wire_man_inf_w_operation_r1_w_range752w(0) <= operation_r1_w(20);
	wire_man_inf_w_operation_r1_w_range754w(0) <= operation_r1_w(21);
	wire_man_inf_w_operation_r1_w_range702w(0) <= operation_r1_w(2);
	wire_man_inf_w_operation_r1_w_range708w(0) <= operation_r1_w(4);
	wire_man_inf_w_operation_r1_w_range710w(0) <= operation_r1_w(5);
	wire_man_inf_w_operation_r1_w_range713w(0) <= operation_r1_w(6);
	wire_man_inf_w_operation_r1_w_range719w(0) <= operation_r1_w(8);
	wire_man_inf_w_operation_r1_w_range721w(0) <= operation_r1_w(9);
	wire_man_inf_w_operation_r2_w_range768w(0) <= operation_r2_w(0);
	wire_man_inf_w_operation_r2_w_range771w(0) <= operation_r2_w(1);
	wire_man_inf_w_operation_r2_w_range774w(0) <= operation_r2_w(2);
	wire_man_inf_w_operation_r2_w_range780w(0) <= operation_r2_w(4);
	wire_man_inf_w_operation_r3_w_range788w(0) <= operation_r3_w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe0 <= ( operation_r1_w(22) & operation_r1_w(19) & operation_r1_w(15) & operation_r1_w(11) & operation_r1_w(7) & operation_r1_w(3));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe1 <= ( operation_r2_w(5) & operation_r2_w(3));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN connection_dffe2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN connection_dffe2(0) <= ( operation_r3_w(1));
			END IF;
		END IF;
	END PROCESS;

 END RTL; --prueba1_altfp_log_and_or_a8b


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="ADD" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=39 aclr clken clock dataa datab result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_csa_s0e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (38 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (38 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (38 DOWNTO 0)
	 ); 
 END prueba1_altfp_log_csa_s0e;

 ARCHITECTURE RTL OF prueba1_altfp_log_csa_s0e IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout803w804w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout802w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout803w804w805w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper0_result	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout803w804w805w & wire_csa_lower_result);
	loop80 : FOR i IN 0 TO 18 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout803w804w(i) <= wire_csa_lower_w_lg_cout803w(0) AND wire_csa_upper0_result(i);
	END GENERATE loop80;
	loop81 : FOR i IN 0 TO 18 GENERATE 
		wire_csa_lower_w_lg_cout802w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop81;
	wire_csa_lower_w_lg_cout803w(0) <= NOT wire_csa_lower_cout;
	loop82 : FOR i IN 0 TO 18 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout803w804w805w(i) <= wire_csa_lower_w_lg_w_lg_cout803w804w(i) OR wire_csa_lower_w_lg_cout802w(i);
	END GENERATE loop82;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 20
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		cout => wire_csa_lower_cout,
		dataa => dataa(19 DOWNTO 0),
		datab => datab(19 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 19
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clken,
		clock => clock,
		dataa => dataa(38 DOWNTO 20),
		datab => datab(38 DOWNTO 20),
		result => wire_csa_upper0_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 19
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_vcc,
		clken => clken,
		clock => clock,
		dataa => dataa(38 DOWNTO 20),
		datab => datab(38 DOWNTO 20),
		result => wire_csa_upper1_result
	  );

 END RTL; --prueba1_altfp_log_csa_s0e


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="ADD" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=31 aclr clken clock dataa datab result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_csa_k0e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (30 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (30 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (30 DOWNTO 0)
	 ); 
 END prueba1_altfp_log_csa_k0e;

 ARCHITECTURE RTL OF prueba1_altfp_log_csa_k0e IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout814w815w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout813w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout814w815w816w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper0_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout814w815w816w & wire_csa_lower_result);
	loop83 : FOR i IN 0 TO 14 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout814w815w(i) <= wire_csa_lower_w_lg_cout814w(0) AND wire_csa_upper0_result(i);
	END GENERATE loop83;
	loop84 : FOR i IN 0 TO 14 GENERATE 
		wire_csa_lower_w_lg_cout813w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop84;
	wire_csa_lower_w_lg_cout814w(0) <= NOT wire_csa_lower_cout;
	loop85 : FOR i IN 0 TO 14 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout814w815w816w(i) <= wire_csa_lower_w_lg_w_lg_cout814w815w(i) OR wire_csa_lower_w_lg_cout813w(i);
	END GENERATE loop85;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 16
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		cout => wire_csa_lower_cout,
		dataa => dataa(15 DOWNTO 0),
		datab => datab(15 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 15
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clken,
		clock => clock,
		dataa => dataa(30 DOWNTO 16),
		datab => datab(30 DOWNTO 16),
		result => wire_csa_upper0_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 15
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_vcc,
		clken => clken,
		clock => clock,
		dataa => dataa(30 DOWNTO 16),
		datab => datab(30 DOWNTO 16),
		result => wire_csa_upper1_result
	  );

 END RTL; --prueba1_altfp_log_csa_k0e


--altfp_log_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=8 dataa datab result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_csa_0nc IS 
	 PORT 
	 ( 
		 dataa	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0)
	 ); 
 END prueba1_altfp_log_csa_0nc;

 ARCHITECTURE RTL OF prueba1_altfp_log_csa_0nc IS

	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub1_result;
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		dataa => dataa,
		datab => datab,
		result => wire_add_sub1_result
	  );

 END RTL; --prueba1_altfp_log_csa_0nc


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=12 dataa datab result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_csa_d4b IS 
	 PORT 
	 ( 
		 dataa	:	IN  STD_LOGIC_VECTOR (11 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (11 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (11 DOWNTO 0)
	 ); 
 END prueba1_altfp_log_csa_d4b;

 ARCHITECTURE RTL OF prueba1_altfp_log_csa_d4b IS

	 SIGNAL  wire_add_sub2_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub2_result;
	add_sub2 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 12
	  )
	  PORT MAP ( 
		dataa => dataa,
		datab => datab,
		result => wire_add_sub2_result
	  );

 END RTL; --prueba1_altfp_log_csa_d4b


--altfp_log_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=6 dataa datab result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_csa_umc IS 
	 PORT 
	 ( 
		 dataa	:	IN  STD_LOGIC_VECTOR (5 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (5 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0)
	 ); 
 END prueba1_altfp_log_csa_umc;

 ARCHITECTURE RTL OF prueba1_altfp_log_csa_umc IS

	 SIGNAL  wire_add_sub3_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub3_result;
	add_sub3 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		dataa => dataa,
		datab => datab,
		result => wire_add_sub3_result
	  );

 END RTL; --prueba1_altfp_log_csa_umc


--altfp_log_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=26 aclr clken clock dataa datab result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_csa_nlf IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (25 DOWNTO 0)
	 ); 
 END prueba1_altfp_log_csa_nlf;

 ARCHITECTURE RTL OF prueba1_altfp_log_csa_nlf IS

	 SIGNAL  wire_add_sub4_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub4_result;
	add_sub4 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 26
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => dataa,
		datab => datab,
		result => wire_add_sub4_result
	  );

 END RTL; --prueba1_altfp_log_csa_nlf


--altfp_log_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_PIPELINE=2 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=8 aclr clken clock dataa datab result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_csa_8kf IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0)
	 ); 
 END prueba1_altfp_log_csa_8kf;

 ARCHITECTURE RTL OF prueba1_altfp_log_csa_8kf IS

	 SIGNAL  wire_add_sub5_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub5_result;
	add_sub5 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 2,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => dataa,
		datab => datab,
		result => wire_add_sub5_result
	  );

 END RTL; --prueba1_altfp_log_csa_8kf


--altfp_log_rr_block CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" WIDTH_ALMOSTLOG=39 WIDTH_Y0=25 WIDTH_Z=26 a0_in aclr almostlog clk_en clock y0_in z
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="ADD" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=29 aclr clken clock dataa datab result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_csa_r0e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (28 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (28 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (28 DOWNTO 0)
	 ); 
 END prueba1_altfp_log_csa_r0e;

 ARCHITECTURE RTL OF prueba1_altfp_log_csa_r0e IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout1203w1204w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1202w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout1203w1204w1205w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper0_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout1203w1204w1205w & wire_csa_lower_result);
	loop86 : FOR i IN 0 TO 13 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout1203w1204w(i) <= wire_csa_lower_w_lg_cout1203w(0) AND wire_csa_upper0_result(i);
	END GENERATE loop86;
	loop87 : FOR i IN 0 TO 13 GENERATE 
		wire_csa_lower_w_lg_cout1202w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop87;
	wire_csa_lower_w_lg_cout1203w(0) <= NOT wire_csa_lower_cout;
	loop88 : FOR i IN 0 TO 13 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout1203w1204w1205w(i) <= wire_csa_lower_w_lg_w_lg_cout1203w1204w(i) OR wire_csa_lower_w_lg_cout1202w(i);
	END GENERATE loop88;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 15
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		cout => wire_csa_lower_cout,
		dataa => dataa(14 DOWNTO 0),
		datab => datab(14 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 14
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clken,
		clock => clock,
		dataa => dataa(28 DOWNTO 15),
		datab => datab(28 DOWNTO 15),
		result => wire_csa_upper0_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 14
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_vcc,
		clken => clken,
		clock => clock,
		dataa => dataa(28 DOWNTO 15),
		datab => datab(28 DOWNTO 15),
		result => wire_csa_upper1_result
	  );

 END RTL; --prueba1_altfp_log_csa_r0e


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="ADD" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=26 aclr clken clock dataa datab result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_csa_o0e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (25 DOWNTO 0)
	 ); 
 END prueba1_altfp_log_csa_o0e;

 ARCHITECTURE RTL OF prueba1_altfp_log_csa_o0e IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout1214w1215w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1213w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout1214w1215w1216w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper0_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout1214w1215w1216w & wire_csa_lower_result);
	loop89 : FOR i IN 0 TO 12 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout1214w1215w(i) <= wire_csa_lower_w_lg_cout1214w(0) AND wire_csa_upper0_result(i);
	END GENERATE loop89;
	loop90 : FOR i IN 0 TO 12 GENERATE 
		wire_csa_lower_w_lg_cout1213w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop90;
	wire_csa_lower_w_lg_cout1214w(0) <= NOT wire_csa_lower_cout;
	loop91 : FOR i IN 0 TO 12 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout1214w1215w1216w(i) <= wire_csa_lower_w_lg_w_lg_cout1214w1215w(i) OR wire_csa_lower_w_lg_cout1213w(i);
	END GENERATE loop91;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		cout => wire_csa_lower_cout,
		dataa => dataa(12 DOWNTO 0),
		datab => datab(12 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clken,
		clock => clock,
		dataa => dataa(25 DOWNTO 13),
		datab => datab(25 DOWNTO 13),
		result => wire_csa_upper0_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_vcc,
		clken => clken,
		clock => clock,
		dataa => dataa(25 DOWNTO 13),
		datab => datab(25 DOWNTO 13),
		result => wire_csa_upper1_result
	  );

 END RTL; --prueba1_altfp_log_csa_o0e


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=31 aclr clken clock dataa datab result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_csa_l1e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (30 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (30 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (30 DOWNTO 0)
	 ); 
 END prueba1_altfp_log_csa_l1e;

 ARCHITECTURE RTL OF prueba1_altfp_log_csa_l1e IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout1225w1226w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1224w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout1225w1226w1227w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper0_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout1225w1226w1227w & wire_csa_lower_result);
	loop92 : FOR i IN 0 TO 14 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout1225w1226w(i) <= wire_csa_lower_w_lg_cout1225w(0) AND wire_csa_upper0_result(i);
	END GENERATE loop92;
	loop93 : FOR i IN 0 TO 14 GENERATE 
		wire_csa_lower_w_lg_cout1224w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop93;
	wire_csa_lower_w_lg_cout1225w(0) <= NOT wire_csa_lower_cout;
	loop94 : FOR i IN 0 TO 14 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout1225w1226w1227w(i) <= wire_csa_lower_w_lg_w_lg_cout1225w1226w(i) OR wire_csa_lower_w_lg_cout1224w(i);
	END GENERATE loop94;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 16
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		cout => wire_csa_lower_cout,
		dataa => dataa(15 DOWNTO 0),
		datab => datab(15 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 15
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clken,
		clock => clock,
		dataa => dataa(30 DOWNTO 16),
		datab => datab(30 DOWNTO 16),
		result => wire_csa_upper0_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 15
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_vcc,
		clken => clken,
		clock => clock,
		dataa => dataa(30 DOWNTO 16),
		datab => datab(30 DOWNTO 16),
		result => wire_csa_upper1_result
	  );

 END RTL; --prueba1_altfp_log_csa_l1e


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=29 aclr clken clock dataa datab result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_csa_s1e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (28 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (28 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (28 DOWNTO 0)
	 ); 
 END prueba1_altfp_log_csa_s1e;

 ARCHITECTURE RTL OF prueba1_altfp_log_csa_s1e IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout1236w1237w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1235w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout1236w1237w1238w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper0_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout1236w1237w1238w & wire_csa_lower_result);
	loop95 : FOR i IN 0 TO 13 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout1236w1237w(i) <= wire_csa_lower_w_lg_cout1236w(0) AND wire_csa_upper0_result(i);
	END GENERATE loop95;
	loop96 : FOR i IN 0 TO 13 GENERATE 
		wire_csa_lower_w_lg_cout1235w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop96;
	wire_csa_lower_w_lg_cout1236w(0) <= NOT wire_csa_lower_cout;
	loop97 : FOR i IN 0 TO 13 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout1236w1237w1238w(i) <= wire_csa_lower_w_lg_w_lg_cout1236w1237w(i) OR wire_csa_lower_w_lg_cout1235w(i);
	END GENERATE loop97;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 15
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		cout => wire_csa_lower_cout,
		dataa => dataa(14 DOWNTO 0),
		datab => datab(14 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 14
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clken,
		clock => clock,
		dataa => dataa(28 DOWNTO 15),
		datab => datab(28 DOWNTO 15),
		result => wire_csa_upper0_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 14
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_vcc,
		clken => clken,
		clock => clock,
		dataa => dataa(28 DOWNTO 15),
		datab => datab(28 DOWNTO 15),
		result => wire_csa_upper1_result
	  );

 END RTL; --prueba1_altfp_log_csa_s1e


--altfp_log_csa CBX_AUTO_BLACKBOX="ALL" LPM_DIRECTION="SUB" LPM_PIPELINE=1 LPM_REPRESENTATION="UNSIGNED" LPM_WIDTH=26 aclr clken clock dataa datab result
--VERSION_BEGIN 15.1 cbx_altbarrel_shift 2015:10:21:18:09:22:SJ cbx_altfp_log 2015:10:21:18:09:22:SJ cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_altsquare 2015:10:21:18:09:23:SJ cbx_cycloneii 2015:10:21:18:09:23:SJ cbx_lpm_add_sub 2015:10:21:18:09:23:SJ cbx_lpm_compare 2015:10:21:18:09:23:SJ cbx_lpm_mult 2015:10:21:18:09:23:SJ cbx_lpm_mux 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ cbx_nadder 2015:10:21:18:09:23:SJ cbx_padd 2015:10:21:18:09:23:SJ cbx_stratix 2015:10:21:18:09:23:SJ cbx_stratixii 2015:10:21:18:09:23:SJ cbx_util_mgl 2015:10:21:18:09:23:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_csa_p1e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (25 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (25 DOWNTO 0)
	 ); 
 END prueba1_altfp_log_csa_p1e;

 ARCHITECTURE RTL OF prueba1_altfp_log_csa_p1e IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout1247w1248w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1246w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout1247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout1247w1248w1249w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper0_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout1247w1248w1249w & wire_csa_lower_result);
	loop98 : FOR i IN 0 TO 12 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout1247w1248w(i) <= wire_csa_lower_w_lg_cout1247w(0) AND wire_csa_upper0_result(i);
	END GENERATE loop98;
	loop99 : FOR i IN 0 TO 12 GENERATE 
		wire_csa_lower_w_lg_cout1246w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop99;
	wire_csa_lower_w_lg_cout1247w(0) <= NOT wire_csa_lower_cout;
	loop100 : FOR i IN 0 TO 12 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout1247w1248w1249w(i) <= wire_csa_lower_w_lg_w_lg_cout1247w1248w(i) OR wire_csa_lower_w_lg_cout1246w(i);
	END GENERATE loop100;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		cout => wire_csa_lower_cout,
		dataa => dataa(12 DOWNTO 0),
		datab => datab(12 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper0 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_gnd,
		clken => clken,
		clock => clock,
		dataa => dataa(25 DOWNTO 13),
		datab => datab(25 DOWNTO 13),
		result => wire_csa_upper0_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aclr => aclr,
		cin => wire_vcc,
		clken => clken,
		clock => clock,
		dataa => dataa(25 DOWNTO 13),
		datab => datab(25 DOWNTO 13),
		result => wire_csa_upper1_result
	  );

 END RTL; --prueba1_altfp_log_csa_p1e

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_add_sub 27 lpm_mult 4 lpm_mux 5 reg 531 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_range_reduction_c2e IS 
	 PORT 
	 ( 
		 a0_in	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 aclr	:	IN  STD_LOGIC := '0';
		 almostlog	:	OUT  STD_LOGIC_VECTOR (38 DOWNTO 0);
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC;
		 y0_in	:	IN  STD_LOGIC_VECTOR (24 DOWNTO 0);
		 z	:	OUT  STD_LOGIC_VECTOR (25 DOWNTO 0)
	 ); 
 END prueba1_range_reduction_c2e;

 ARCHITECTURE RTL OF prueba1_range_reduction_c2e IS

	 SIGNAL  wire_add0_1_datab	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add0_1_result	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add0_2_datab	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add0_2_result	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add0_3_datab	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add0_3_result	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add1_1_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add1_2_result	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_add1_3_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_sub1_1_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_sub1_2_result	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_sub1_3_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL	 A_pipe0_reg0	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 A_pipe0_reg1	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 A_pipe0_reg2	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 A_wire1_reg0	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 A_wire2_reg0	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 A_wire3_reg0	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 B_wire1_reg0	:	STD_LOGIC_VECTOR(20 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 B_wire2_reg0	:	STD_LOGIC_VECTOR(26 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 B_wire3_reg0	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 P_pipe0_reg0	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 P_pipe1_reg0	:	STD_LOGIC_VECTOR(28 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 P_pipe2_reg0	:	STD_LOGIC_VECTOR(28 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 P_pipe3_reg0	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 S_pipe22_reg0	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 S_pipe23_reg0	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 S_pipe24_reg0	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 S_wire1_reg0	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 S_wire2_reg0	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 S_wire3_reg0	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Z_wire1_reg0	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Z_wire2_reg0	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Z_wire3_reg0	:	STD_LOGIC_VECTOR(28 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_mult0_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_mult1_result	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_mult2_result	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_mult3_result	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_InvTable0_data	:	STD_LOGIC_VECTOR (191 DOWNTO 0);
	 SIGNAL  wire_InvTable0_data_2d	:	STD_LOGIC_2D(31 DOWNTO 0, 5 DOWNTO 0);
	 SIGNAL  wire_InvTable0_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_LogTable0_data	:	STD_LOGIC_VECTOR (1247 DOWNTO 0);
	 SIGNAL  wire_LogTable0_data_2d	:	STD_LOGIC_2D(31 DOWNTO 0, 38 DOWNTO 0);
	 SIGNAL  wire_LogTable0_result	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_LogTable1_data	:	STD_LOGIC_VECTOR (559 DOWNTO 0);
	 SIGNAL  wire_LogTable1_data_2d	:	STD_LOGIC_2D(15 DOWNTO 0, 34 DOWNTO 0);
	 SIGNAL  wire_LogTable1_result	:	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  wire_LogTable2_data	:	STD_LOGIC_VECTOR (511 DOWNTO 0);
	 SIGNAL  wire_LogTable2_data_2d	:	STD_LOGIC_2D(15 DOWNTO 0, 31 DOWNTO 0);
	 SIGNAL  wire_LogTable2_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_LogTable3_data	:	STD_LOGIC_VECTOR (463 DOWNTO 0);
	 SIGNAL  wire_LogTable3_data_2d	:	STD_LOGIC_2D(15 DOWNTO 0, 28 DOWNTO 0);
	 SIGNAL  wire_LogTable3_result	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A1_is_not_zero_range1009w1027w1028w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_all_zero2_range1099w1103w1107w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_all_zero3_range1176w1180w1184w	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_pipe11_range1004w1007w1008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1088w1089w1090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1092w1093w1094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1096w1097w1098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1165w1166w1167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1169w1170w1171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1173w1174w1175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A1_is_all_zero_range1006w1030w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A1_is_not_zero_range1009w1026w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A1_is_not_zero_range1009w1027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_all_zero2_range1099w1103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_all_zero3_range1176w1180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe11_range1004w1007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe12_range1084w1085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe12_range1088w1089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe12_range1092w1093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe12_range1096w1097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe13_range1161w1162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe13_range1165w1166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe13_range1169w1170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe13_range1173w1174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w1029w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe11_range994w995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe11_range994w997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe11_range999w1000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe11_range999w1002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_lg_w_A_pipe11_range1004w1005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  A1_is_all_zero :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A1_is_not_zero :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_all_zero2 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_all_zero3 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_pipe0 :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  A_pipe11 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_pipe12 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_pipe13 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_wire0 :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  A_wire1 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_wire2 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  A_wire3 :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  B_pad_wire1 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  B_pad_wire2 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  B_pad_wire3 :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  B_pipe1 :	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  B_pipe2 :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  B_pipe3 :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  B_wire1 :	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  B_wire2 :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  B_wire3 :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  epsZ_pad_wire1 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  epsZ_pad_wire2 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  epsZ_pad_wire3 :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  epsZ_wire1 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  epsZ_wire2 :	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  epsZ_wire3 :	STD_LOGIC_VECTOR (40 DOWNTO 0);
	 SIGNAL  InvA0 :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  L_wire0 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  L_wire1 :	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  L_wire2 :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  L_wire3 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  mux0_data0 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  mux0_data1 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  P_pad_wire1 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  P_pad_wire2 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  P_pad_wire3 :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  P_pipe0 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  P_pipe1 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  P_pipe2 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  P_pipe3 :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  P_wire0 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  P_wire1 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  P_wire2 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  P_wire3 :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  S_pipe11 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_pipe12 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_pipe13 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_pipe22 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_pipe23 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_pipe24 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_wire1 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_wire2 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_wire3 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  S_wire4 :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  Z_pipe1 :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Z_pipe2 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  Z_pipe3 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  Z_wire1 :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Z_wire2 :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  Z_wire3 :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  Z_wire4 :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  ZM_wire1 :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  ZM_wire2 :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  ZM_wire3 :	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_all_zero_range990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_all_zero_range996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_all_zero_range1001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_all_zero_range1006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_not_zero_range992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_not_zero_range998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_not_zero_range1003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A1_is_not_zero_range1009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero2_range1086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero2_range1091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero2_range1095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero2_range1099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero3_range1163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero3_range1168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero3_range1172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_all_zero3_range1176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe11_range994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe11_range999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe11_range1004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe12_range1084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe12_range1088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe12_range1092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe12_range1096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe13_range1161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe13_range1165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe13_range1169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_range_reduction_w_A_pipe13_range1173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  prueba1_altfp_log_csa_s0e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(38 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(38 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(38 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_csa_k0e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(30 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(30 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(30 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_csa_r0e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(28 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(28 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(28 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_csa_o0e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(25 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_csa_l1e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(30 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(30 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(30 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_csa_s1e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(28 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(28 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(28 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_csa_p1e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(25 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop101 : FOR i IN 0 TO 30 GENERATE 
		wire_range_reduction_w_lg_w_lg_w_A1_is_not_zero_range1009w1027w1028w(i) <= wire_range_reduction_w_lg_w_A1_is_not_zero_range1009w1027w(0) AND mux0_data0(i);
	END GENERATE loop101;
	loop102 : FOR i IN 0 TO 30 GENERATE 
		wire_range_reduction_w_lg_w_lg_w_A_all_zero2_range1099w1103w1107w(i) <= wire_range_reduction_w_lg_w_A_all_zero2_range1099w1103w(0) AND Z_pipe2(i);
	END GENERATE loop102;
	loop103 : FOR i IN 0 TO 28 GENERATE 
		wire_range_reduction_w_lg_w_lg_w_A_all_zero3_range1176w1180w1184w(i) <= wire_range_reduction_w_lg_w_A_all_zero3_range1176w1180w(0) AND Z_pipe3(i);
	END GENERATE loop103;
	wire_range_reduction_w_lg_w_lg_w_A_pipe11_range1004w1007w1008w(0) <= wire_range_reduction_w_lg_w_A_pipe11_range1004w1007w(0) AND wire_range_reduction_w_A1_is_not_zero_range1003w(0);
	wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1088w1089w1090w(0) <= wire_range_reduction_w_lg_w_A_pipe12_range1088w1089w(0) AND wire_range_reduction_w_A_all_zero2_range1086w(0);
	wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1092w1093w1094w(0) <= wire_range_reduction_w_lg_w_A_pipe12_range1092w1093w(0) AND wire_range_reduction_w_A_all_zero2_range1091w(0);
	wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1096w1097w1098w(0) <= wire_range_reduction_w_lg_w_A_pipe12_range1096w1097w(0) AND wire_range_reduction_w_A_all_zero2_range1095w(0);
	wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1165w1166w1167w(0) <= wire_range_reduction_w_lg_w_A_pipe13_range1165w1166w(0) AND wire_range_reduction_w_A_all_zero3_range1163w(0);
	wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1169w1170w1171w(0) <= wire_range_reduction_w_lg_w_A_pipe13_range1169w1170w(0) AND wire_range_reduction_w_A_all_zero3_range1168w(0);
	wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1173w1174w1175w(0) <= wire_range_reduction_w_lg_w_A_pipe13_range1173w1174w(0) AND wire_range_reduction_w_A_all_zero3_range1172w(0);
	loop104 : FOR i IN 0 TO 30 GENERATE 
		wire_range_reduction_w_lg_w_A1_is_all_zero_range1006w1030w(i) <= wire_range_reduction_w_A1_is_all_zero_range1006w(0) AND wire_range_reduction_w1029w(i);
	END GENERATE loop104;
	loop105 : FOR i IN 0 TO 30 GENERATE 
		wire_range_reduction_w_lg_w_A1_is_not_zero_range1009w1026w(i) <= wire_range_reduction_w_A1_is_not_zero_range1009w(0) AND mux0_data1(i);
	END GENERATE loop105;
	wire_range_reduction_w_lg_w_A1_is_not_zero_range1009w1027w(0) <= NOT wire_range_reduction_w_A1_is_not_zero_range1009w(0);
	wire_range_reduction_w_lg_w_A_all_zero2_range1099w1103w(0) <= NOT wire_range_reduction_w_A_all_zero2_range1099w(0);
	wire_range_reduction_w_lg_w_A_all_zero3_range1176w1180w(0) <= NOT wire_range_reduction_w_A_all_zero3_range1176w(0);
	wire_range_reduction_w_lg_w_A_pipe11_range1004w1007w(0) <= NOT wire_range_reduction_w_A_pipe11_range1004w(0);
	wire_range_reduction_w_lg_w_A_pipe12_range1084w1085w(0) <= NOT wire_range_reduction_w_A_pipe12_range1084w(0);
	wire_range_reduction_w_lg_w_A_pipe12_range1088w1089w(0) <= NOT wire_range_reduction_w_A_pipe12_range1088w(0);
	wire_range_reduction_w_lg_w_A_pipe12_range1092w1093w(0) <= NOT wire_range_reduction_w_A_pipe12_range1092w(0);
	wire_range_reduction_w_lg_w_A_pipe12_range1096w1097w(0) <= NOT wire_range_reduction_w_A_pipe12_range1096w(0);
	wire_range_reduction_w_lg_w_A_pipe13_range1161w1162w(0) <= NOT wire_range_reduction_w_A_pipe13_range1161w(0);
	wire_range_reduction_w_lg_w_A_pipe13_range1165w1166w(0) <= NOT wire_range_reduction_w_A_pipe13_range1165w(0);
	wire_range_reduction_w_lg_w_A_pipe13_range1169w1170w(0) <= NOT wire_range_reduction_w_A_pipe13_range1169w(0);
	wire_range_reduction_w_lg_w_A_pipe13_range1173w1174w(0) <= NOT wire_range_reduction_w_A_pipe13_range1173w(0);
	loop106 : FOR i IN 0 TO 30 GENERATE 
		wire_range_reduction_w1029w(i) <= wire_range_reduction_w_lg_w_lg_w_A1_is_not_zero_range1009w1027w1028w(i) OR wire_range_reduction_w_lg_w_A1_is_not_zero_range1009w1026w(i);
	END GENERATE loop106;
	wire_range_reduction_w_lg_w_A_pipe11_range994w995w(0) <= wire_range_reduction_w_A_pipe11_range994w(0) OR wire_range_reduction_w_A1_is_all_zero_range990w(0);
	wire_range_reduction_w_lg_w_A_pipe11_range994w997w(0) <= wire_range_reduction_w_A_pipe11_range994w(0) OR wire_range_reduction_w_A1_is_not_zero_range992w(0);
	wire_range_reduction_w_lg_w_A_pipe11_range999w1000w(0) <= wire_range_reduction_w_A_pipe11_range999w(0) OR wire_range_reduction_w_A1_is_all_zero_range996w(0);
	wire_range_reduction_w_lg_w_A_pipe11_range999w1002w(0) <= wire_range_reduction_w_A_pipe11_range999w(0) OR wire_range_reduction_w_A1_is_not_zero_range998w(0);
	wire_range_reduction_w_lg_w_A_pipe11_range1004w1005w(0) <= wire_range_reduction_w_A_pipe11_range1004w(0) OR wire_range_reduction_w_A1_is_all_zero_range1001w(0);
	A1_is_all_zero <= ( wire_range_reduction_w_lg_w_A_pipe11_range1004w1005w & wire_range_reduction_w_lg_w_A_pipe11_range999w1000w & wire_range_reduction_w_lg_w_A_pipe11_range994w995w & A_pipe11(0));
	A1_is_not_zero <= ( wire_range_reduction_w_lg_w_lg_w_A_pipe11_range1004w1007w1008w & wire_range_reduction_w_lg_w_A_pipe11_range999w1002w & wire_range_reduction_w_lg_w_A_pipe11_range994w997w & A_pipe11(0));
	A_all_zero2 <= ( wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1096w1097w1098w & wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1092w1093w1094w & wire_range_reduction_w_lg_w_lg_w_A_pipe12_range1088w1089w1090w & wire_range_reduction_w_lg_w_A_pipe12_range1084w1085w);
	A_all_zero3 <= ( wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1173w1174w1175w & wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1169w1170w1171w & wire_range_reduction_w_lg_w_lg_w_A_pipe13_range1165w1166w1167w & wire_range_reduction_w_lg_w_A_pipe13_range1161w1162w);
	A_pipe0 <= a0_in;
	A_pipe11 <= A_wire1_reg0;
	A_pipe12 <= A_wire2_reg0;
	A_pipe13 <= A_wire3_reg0;
	A_wire0 <= A_pipe0_reg2;
	A_wire1 <= Z_wire1(24 DOWNTO 21);
	A_wire2 <= Z_wire2(30 DOWNTO 27);
	A_wire3 <= Z_wire3(28 DOWNTO 25);
	almostlog <= S_wire4;
	B_pad_wire1 <= ( "0" & B_pipe1 & "000000000");
	B_pad_wire2 <= ( "0" & B_pipe2 & "0");
	B_pad_wire3 <= ( "0" & B_pipe3);
	B_pipe1 <= B_wire1_reg0;
	B_pipe2 <= B_wire2_reg0;
	B_pipe3 <= B_wire3_reg0;
	B_wire1 <= Z_wire1(20 DOWNTO 0);
	B_wire2 <= Z_wire2(26 DOWNTO 0);
	B_wire3 <= Z_wire3(24 DOWNTO 0);
	epsZ_pad_wire1 <= epsZ_wire1(30 DOWNTO 0);
	epsZ_pad_wire2 <= epsZ_wire2(39 DOWNTO 11);
	epsZ_pad_wire3 <= epsZ_wire3(40 DOWNTO 15);
	epsZ_wire1 <= wire_range_reduction_w_lg_w_A1_is_all_zero_range1006w1030w;
	epsZ_wire2 <= ( "0" & wire_range_reduction_w_lg_w_A_all_zero2_range1099w1103w & "0000000" & wire_range_reduction_w_lg_w_lg_w_A_all_zero2_range1099w1103w1107w);
	epsZ_wire3 <= ( "0" & wire_range_reduction_w_lg_w_A_all_zero3_range1176w1180w & "0000000000" & wire_range_reduction_w_lg_w_lg_w_A_all_zero3_range1176w1180w1184w);
	InvA0 <= wire_InvTable0_result;
	L_wire0 <= wire_LogTable0_result;
	L_wire1 <= wire_LogTable1_result;
	L_wire2 <= wire_LogTable2_result;
	L_wire3 <= wire_LogTable3_result;
	mux0_data0 <= ( "1" & "0000" & Z_pipe1 & "0");
	mux0_data1 <= ( "0" & "1" & "0000" & Z_pipe1);
	P_pad_wire1 <= ( "0" & P_wire1 & "0");
	P_pad_wire2 <= ( "0000" & P_wire2(28 DOWNTO 4));
	P_pad_wire3 <= ( "0000000" & P_wire3(22 DOWNTO 4));
	P_pipe0 <= wire_mult0_result;
	P_pipe1 <= wire_mult1_result;
	P_pipe2 <= wire_mult2_result;
	P_pipe3 <= wire_mult3_result;
	P_wire0 <= P_pipe0_reg0;
	P_wire1 <= P_pipe1_reg0;
	P_wire2 <= P_pipe2_reg0;
	P_wire3 <= P_pipe3_reg0;
	S_pipe11 <= S_wire1_reg0;
	S_pipe12 <= S_wire2_reg0;
	S_pipe13 <= S_wire3_reg0;
	S_pipe22 <= wire_add0_1_result;
	S_pipe23 <= wire_add0_2_result;
	S_pipe24 <= wire_add0_3_result;
	S_wire1 <= L_wire0;
	S_wire2 <= S_pipe22_reg0;
	S_wire3 <= S_pipe23_reg0;
	S_wire4 <= S_pipe24_reg0;
	z <= Z_wire4;
	Z_pipe1 <= Z_wire1_reg0;
	Z_pipe2 <= Z_wire2_reg0;
	Z_pipe3 <= Z_wire3_reg0;
	Z_wire1 <= P_wire0(24 DOWNTO 0);
	Z_wire2 <= wire_sub1_1_result;
	Z_wire3 <= wire_sub1_2_result;
	Z_wire4 <= wire_sub1_3_result;
	ZM_wire1 <= Z_wire1;
	ZM_wire2 <= Z_wire2(30 DOWNTO 6);
	ZM_wire3 <= Z_wire3(28 DOWNTO 10);
	wire_range_reduction_w_A1_is_all_zero_range990w(0) <= A1_is_all_zero(0);
	wire_range_reduction_w_A1_is_all_zero_range996w(0) <= A1_is_all_zero(1);
	wire_range_reduction_w_A1_is_all_zero_range1001w(0) <= A1_is_all_zero(2);
	wire_range_reduction_w_A1_is_all_zero_range1006w(0) <= A1_is_all_zero(3);
	wire_range_reduction_w_A1_is_not_zero_range992w(0) <= A1_is_not_zero(0);
	wire_range_reduction_w_A1_is_not_zero_range998w(0) <= A1_is_not_zero(1);
	wire_range_reduction_w_A1_is_not_zero_range1003w(0) <= A1_is_not_zero(2);
	wire_range_reduction_w_A1_is_not_zero_range1009w(0) <= A1_is_not_zero(3);
	wire_range_reduction_w_A_all_zero2_range1086w(0) <= A_all_zero2(0);
	wire_range_reduction_w_A_all_zero2_range1091w(0) <= A_all_zero2(1);
	wire_range_reduction_w_A_all_zero2_range1095w(0) <= A_all_zero2(2);
	wire_range_reduction_w_A_all_zero2_range1099w(0) <= A_all_zero2(3);
	wire_range_reduction_w_A_all_zero3_range1163w(0) <= A_all_zero3(0);
	wire_range_reduction_w_A_all_zero3_range1168w(0) <= A_all_zero3(1);
	wire_range_reduction_w_A_all_zero3_range1172w(0) <= A_all_zero3(2);
	wire_range_reduction_w_A_all_zero3_range1176w(0) <= A_all_zero3(3);
	wire_range_reduction_w_A_pipe11_range994w(0) <= A_pipe11(1);
	wire_range_reduction_w_A_pipe11_range999w(0) <= A_pipe11(2);
	wire_range_reduction_w_A_pipe11_range1004w(0) <= A_pipe11(3);
	wire_range_reduction_w_A_pipe12_range1084w(0) <= A_pipe12(0);
	wire_range_reduction_w_A_pipe12_range1088w(0) <= A_pipe12(1);
	wire_range_reduction_w_A_pipe12_range1092w(0) <= A_pipe12(2);
	wire_range_reduction_w_A_pipe12_range1096w(0) <= A_pipe12(3);
	wire_range_reduction_w_A_pipe13_range1161w(0) <= A_pipe13(0);
	wire_range_reduction_w_A_pipe13_range1165w(0) <= A_pipe13(1);
	wire_range_reduction_w_A_pipe13_range1169w(0) <= A_pipe13(2);
	wire_range_reduction_w_A_pipe13_range1173w(0) <= A_pipe13(3);
	wire_add0_1_datab <= ( "0000" & L_wire1);
	add0_1 :  prueba1_altfp_log_csa_s0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => S_pipe11,
		datab => wire_add0_1_datab,
		result => wire_add0_1_result
	  );
	wire_add0_2_datab <= ( "0000000" & L_wire2);
	add0_2 :  prueba1_altfp_log_csa_s0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => S_pipe12,
		datab => wire_add0_2_datab,
		result => wire_add0_2_result
	  );
	wire_add0_3_datab <= ( "0000000000" & L_wire3);
	add0_3 :  prueba1_altfp_log_csa_s0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => S_pipe13,
		datab => wire_add0_3_datab,
		result => wire_add0_3_result
	  );
	add1_1 :  prueba1_altfp_log_csa_k0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => B_pad_wire1,
		datab => epsZ_pad_wire1,
		result => wire_add1_1_result
	  );
	add1_2 :  prueba1_altfp_log_csa_r0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => B_pad_wire2,
		datab => epsZ_pad_wire2,
		result => wire_add1_2_result
	  );
	add1_3 :  prueba1_altfp_log_csa_o0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => B_pad_wire3,
		datab => epsZ_pad_wire3,
		result => wire_add1_3_result
	  );
	sub1_1 :  prueba1_altfp_log_csa_l1e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_add1_1_result,
		datab => P_pad_wire1,
		result => wire_sub1_1_result
	  );
	sub1_2 :  prueba1_altfp_log_csa_s1e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_add1_2_result,
		datab => P_pad_wire2,
		result => wire_sub1_2_result
	  );
	sub1_3 :  prueba1_altfp_log_csa_p1e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_add1_3_result,
		datab => P_pad_wire3,
		result => wire_sub1_3_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN A_pipe0_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN A_pipe0_reg0 <= A_pipe0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN A_pipe0_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN A_pipe0_reg1 <= A_pipe0_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN A_pipe0_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN A_pipe0_reg2 <= A_pipe0_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN A_wire1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN A_wire1_reg0 <= A_wire1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN A_wire2_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN A_wire2_reg0 <= A_wire2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN A_wire3_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN A_wire3_reg0 <= A_wire3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN B_wire1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN B_wire1_reg0 <= B_wire1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN B_wire2_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN B_wire2_reg0 <= B_wire2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN B_wire3_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN B_wire3_reg0 <= B_wire3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN P_pipe0_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN P_pipe0_reg0 <= P_pipe0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN P_pipe1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN P_pipe1_reg0 <= P_pipe1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN P_pipe2_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN P_pipe2_reg0 <= P_pipe2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN P_pipe3_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN P_pipe3_reg0 <= P_pipe3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN S_pipe22_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN S_pipe22_reg0 <= S_pipe22;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN S_pipe23_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN S_pipe23_reg0 <= S_pipe23;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN S_pipe24_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN S_pipe24_reg0 <= S_pipe24;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN S_wire1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN S_wire1_reg0 <= S_wire1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN S_wire2_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN S_wire2_reg0 <= S_wire2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN S_wire3_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN S_wire3_reg0 <= S_wire3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Z_wire1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Z_wire1_reg0 <= Z_wire1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Z_wire2_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Z_wire2_reg0 <= Z_wire2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Z_wire3_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Z_wire3_reg0 <= Z_wire3;
			END IF;
		END IF;
	END PROCESS;
	mult0 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 2,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 6,
		LPM_WIDTHB => 25,
		LPM_WIDTHP => 31
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => InvA0,
		datab => y0_in,
		result => wire_mult0_result
	  );
	mult1 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 4,
		LPM_WIDTHB => 25,
		LPM_WIDTHP => 29
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => A_wire1,
		datab => ZM_wire1,
		result => wire_mult1_result
	  );
	mult2 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 4,
		LPM_WIDTHB => 25,
		LPM_WIDTHP => 29
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => A_wire2,
		datab => ZM_wire2,
		result => wire_mult2_result
	  );
	mult3 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 4,
		LPM_WIDTHB => 19,
		LPM_WIDTHP => 23
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => A_wire3,
		datab => ZM_wire3,
		result => wire_mult3_result
	  );
	wire_InvTable0_data <= ( "100001" & "100010" & "100010" & "100011" & "100011" & "100100" & "100100" & "100101" & "100110" & "100110" & "100111" & "101000" & "101001" & "101001" & "101010" & "101011" & "010110" & "010111" & "010111" & "011000" & "011000" & "011001" & "011001" & "011010" & "011011" & "011011" & "011100" & "011101" & "011110" & "011111" & "100000" & "100000");
	loop107 : FOR i IN 0 TO 31 GENERATE
		loop108 : FOR j IN 0 TO 5 GENERATE
			wire_InvTable0_data_2d(i, j) <= wire_InvTable0_data(i*6+j);
		END GENERATE loop108;
	END GENERATE loop107;
	InvTable0 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 32,
		LPM_WIDTH => 6,
		LPM_WIDTHS => 5
	  )
	  PORT MAP ( 
		data => wire_InvTable0_data_2d,
		result => wire_InvTable0_result,
		sel => a0_in
	  );
	wire_LogTable0_data <= ( "111110000001111101011001001111000110001" & "111100000111101011100111100111111111100" & "111100000111101011100111100111111111100" & "111010010000111100101101011101010001110" & "111010010000111100101101011101010001110" & "111000011101100011111000100100011101011" & "111000011101100011111000100100011101011" & "110110101101010101011010000011111100001" & "110101000000000110011111000111101011001" & "110101000000000110011111000111101011001" & "110011010101101101001010110001100001100" & "110001101110000000010000011100001100110" & "110000001000110111001111001001010100010" & "110000001000110111001111001001010100010" & "101110100110001010001101010100010101001" & "101101000101110001110101000101000111110" & "010111111110101111101000111011110110000" & "010101001000101010111000000111001110001" & "010101001000101010111000000111001110001" & "010010011010010110001000010001001101001" & "010010011010010110001000010001001101001" & "001111110011001000111000110110010110011" & "001111110011001000111000110110010110011" & "001101010010011111011010011110010001010" & "001010110111111010000000110101101010100" & "001010110111111010000000110101101010100" & "001000100010111100011101000001000100111" & "000110010011001101011110010111010101100" & "000100001000010110011000101101011001111" & "000010000010000010101110110001001111001" & "000000000000000000000000000000000000000" & "000000000000000000000000000000000000000");
	loop109 : FOR i IN 0 TO 31 GENERATE
		loop110 : FOR j IN 0 TO 38 GENERATE
			wire_LogTable0_data_2d(i, j) <= wire_LogTable0_data(i*39+j);
		END GENERATE loop110;
	END GENERATE loop109;
	LogTable0 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 32,
		LPM_WIDTH => 39,
		LPM_WIDTHS => 5
	  )
	  PORT MAP ( 
		data => wire_LogTable0_data_2d,
		result => wire_LogTable0_result,
		sel => A_wire0
	  );
	wire_LogTable1_data <= ( "11100110010110111001111001101110111" & "11010101011101111001011010000111110" & "11000100101001010101000010100100111" & "10110011111001001010011110010110101" & "10100011001101010111011010100001011" & "10010010100101111001100101111100011" & "10000010000010101110110001001111001" & "01110001100011110100101110110000010" & "01101001010101111101010100100011000" & "01011000111101011000010111100001101" & "01001000101000111110110001111111101" & "00111000011000101110011100001001100" & "00101000001100100101001111110010110" & "00011000000100100001001000010100010" & "00001000000000100000000010101010111" & "00000000000000000000000000000000000");
	loop111 : FOR i IN 0 TO 15 GENERATE
		loop112 : FOR j IN 0 TO 34 GENERATE
			wire_LogTable1_data_2d(i, j) <= wire_LogTable1_data(i*35+j);
		END GENERATE loop112;
	END GENERATE loop111;
	LogTable1 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 16,
		LPM_WIDTH => 35,
		LPM_WIDTHS => 4
	  )
	  PORT MAP ( 
		data => wire_LogTable1_data_2d,
		result => wire_LogTable1_result,
		sel => A_pipe11
	  );
	wire_LogTable2_data <= ( "11101000110100110011111101101000" & "11011000101101110000111000001100" & "11001000100111001110001110000010" & "10111000100001001011111101000110" & "10101000011011101010000011010111" & "10011000010110101000011110110010" & "10001000010010000111001101010110" & "01111000001110000110001101000000" & "01101000001010100101011011110000" & "01011000000111100100110111100100" & "01001000000101000100011110011011" & "00111000000011000100001110010011" & "00101000000001100100000101001101" & "00011000000000100100000001001000" & "00001000000000000100000000000010" & "00000000000000000000000000000000");
	loop113 : FOR i IN 0 TO 15 GENERATE
		loop114 : FOR j IN 0 TO 31 GENERATE
			wire_LogTable2_data_2d(i, j) <= wire_LogTable2_data(i*32+j);
		END GENERATE loop114;
	END GENERATE loop113;
	LogTable2 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 16,
		LPM_WIDTH => 32,
		LPM_WIDTHS => 4
	  )
	  PORT MAP ( 
		data => wire_LogTable2_data_2d,
		result => wire_LogTable2_result,
		sel => A_pipe12
	  );
	wire_LogTable3_data <= ( "11101000000110100100101111111" & "11011000000101101100101100110" & "11001000000100111000101010001" & "10111000000100001000100111111" & "10101000000011011100100110000" & "10011000000010110100100100011" & "10001000000010010000100011001" & "01111000000001110000100010001" & "01101000000001010100100001011" & "01011000000000111100100000110" & "01001000000000101000100000011" & "00111000000000011000100000001" & "00101000000000001100100000000" & "00011000000000000100100000000" & "00001000000000000000100000000" & "00000000000000000000000000000");
	loop115 : FOR i IN 0 TO 15 GENERATE
		loop116 : FOR j IN 0 TO 28 GENERATE
			wire_LogTable3_data_2d(i, j) <= wire_LogTable3_data(i*29+j);
		END GENERATE loop116;
	END GENERATE loop115;
	LogTable3 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 16,
		LPM_WIDTH => 29,
		LPM_WIDTHS => 4
	  )
	  PORT MAP ( 
		data => wire_LogTable3_data_2d,
		result => wire_LogTable3_result,
		sel => A_pipe13
	  );

 END RTL; --prueba1_range_reduction_c2e


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" PIPELINE=1 WIDTH=64 WIDTHAD=6 aclr clk_en clock data q
--VERSION_BEGIN 15.1 cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" PIPELINE=0 WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 15.1 cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q
--VERSION_BEGIN 15.1 cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q
--VERSION_BEGIN 15.1 cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q
--VERSION_BEGIN 15.1 cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q
--VERSION_BEGIN 15.1 cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altpriority_encoder_3v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0)
	 ); 
 END prueba1_altpriority_encoder_3v7;

 ARCHITECTURE RTL OF prueba1_altpriority_encoder_3v7 IS

 BEGIN

	q(0) <= ( data(1));

 END RTL; --prueba1_altpriority_encoder_3v7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q zero
--VERSION_BEGIN 15.1 cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altpriority_encoder_3e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END prueba1_altpriority_encoder_3e8;

 ARCHITECTURE RTL OF prueba1_altpriority_encoder_3e8 IS

 BEGIN

	q(0) <= ( data(1));
	zero <= (NOT (data(0) OR data(1)));

 END RTL; --prueba1_altpriority_encoder_3e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altpriority_encoder_6v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0)
	 ); 
 END prueba1_altpriority_encoder_6v7;

 ARCHITECTURE RTL OF prueba1_altpriority_encoder_6v7 IS

	 SIGNAL  wire_altpriority_encoder14_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_w_lg_w_lg_zero1290w1291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_w_lg_zero1292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_w_lg_zero1290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_w_lg_w_lg_zero1292w1293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_zero	:	STD_LOGIC;
	 COMPONENT  prueba1_altpriority_encoder_3v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder15_w_lg_zero1290w & wire_altpriority_encoder15_w_lg_w_lg_zero1292w1293w);
	altpriority_encoder14 :  prueba1_altpriority_encoder_3v7
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder14_q
	  );
	wire_altpriority_encoder15_w_lg_w_lg_zero1290w1291w(0) <= wire_altpriority_encoder15_w_lg_zero1290w(0) AND wire_altpriority_encoder15_q(0);
	wire_altpriority_encoder15_w_lg_zero1292w(0) <= wire_altpriority_encoder15_zero AND wire_altpriority_encoder14_q(0);
	wire_altpriority_encoder15_w_lg_zero1290w(0) <= NOT wire_altpriority_encoder15_zero;
	wire_altpriority_encoder15_w_lg_w_lg_zero1292w1293w(0) <= wire_altpriority_encoder15_w_lg_zero1292w(0) OR wire_altpriority_encoder15_w_lg_w_lg_zero1290w1291w(0);
	altpriority_encoder15 :  prueba1_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder15_q,
		zero => wire_altpriority_encoder15_zero
	  );

 END RTL; --prueba1_altpriority_encoder_6v7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q zero
--VERSION_BEGIN 15.1 cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altpriority_encoder_6e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END prueba1_altpriority_encoder_6e8;

 ARCHITECTURE RTL OF prueba1_altpriority_encoder_6e8 IS

	 SIGNAL  wire_altpriority_encoder16_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder17_w_lg_w_lg_zero1308w1309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_w_lg_zero1310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_w_lg_zero1308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_w_lg_w_lg_zero1310w1311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder17_zero	:	STD_LOGIC;
	 COMPONENT  prueba1_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder17_w_lg_zero1308w & wire_altpriority_encoder17_w_lg_w_lg_zero1310w1311w);
	zero <= (wire_altpriority_encoder16_zero AND wire_altpriority_encoder17_zero);
	altpriority_encoder16 :  prueba1_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder16_q,
		zero => wire_altpriority_encoder16_zero
	  );
	wire_altpriority_encoder17_w_lg_w_lg_zero1308w1309w(0) <= wire_altpriority_encoder17_w_lg_zero1308w(0) AND wire_altpriority_encoder17_q(0);
	wire_altpriority_encoder17_w_lg_zero1310w(0) <= wire_altpriority_encoder17_zero AND wire_altpriority_encoder16_q(0);
	wire_altpriority_encoder17_w_lg_zero1308w(0) <= NOT wire_altpriority_encoder17_zero;
	wire_altpriority_encoder17_w_lg_w_lg_zero1310w1311w(0) <= wire_altpriority_encoder17_w_lg_zero1310w(0) OR wire_altpriority_encoder17_w_lg_w_lg_zero1308w1309w(0);
	altpriority_encoder17 :  prueba1_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder17_q,
		zero => wire_altpriority_encoder17_zero
	  );

 END RTL; --prueba1_altpriority_encoder_6e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altpriority_encoder_bv7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END prueba1_altpriority_encoder_bv7;

 ARCHITECTURE RTL OF prueba1_altpriority_encoder_bv7 IS

	 SIGNAL  wire_altpriority_encoder12_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_w_lg_w_lg_zero1281w1282w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_w_lg_zero1283w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_w_lg_zero1281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_w_lg_w_lg_zero1283w1284w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_zero	:	STD_LOGIC;
	 COMPONENT  prueba1_altpriority_encoder_6v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder13_w_lg_zero1281w & wire_altpriority_encoder13_w_lg_w_lg_zero1283w1284w);
	altpriority_encoder12 :  prueba1_altpriority_encoder_6v7
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder12_q
	  );
	loop117 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder13_w_lg_w_lg_zero1281w1282w(i) <= wire_altpriority_encoder13_w_lg_zero1281w(0) AND wire_altpriority_encoder13_q(i);
	END GENERATE loop117;
	loop118 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder13_w_lg_zero1283w(i) <= wire_altpriority_encoder13_zero AND wire_altpriority_encoder12_q(i);
	END GENERATE loop118;
	wire_altpriority_encoder13_w_lg_zero1281w(0) <= NOT wire_altpriority_encoder13_zero;
	loop119 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder13_w_lg_w_lg_zero1283w1284w(i) <= wire_altpriority_encoder13_w_lg_zero1283w(i) OR wire_altpriority_encoder13_w_lg_w_lg_zero1281w1282w(i);
	END GENERATE loop119;
	altpriority_encoder13 :  prueba1_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder13_q,
		zero => wire_altpriority_encoder13_zero
	  );

 END RTL; --prueba1_altpriority_encoder_bv7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q zero
--VERSION_BEGIN 15.1 cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altpriority_encoder_be8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END prueba1_altpriority_encoder_be8;

 ARCHITECTURE RTL OF prueba1_altpriority_encoder_be8 IS

	 SIGNAL  wire_altpriority_encoder18_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder19_w_lg_w_lg_zero1318w1319w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_w_lg_zero1320w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_w_lg_zero1318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_w_lg_w_lg_zero1320w1321w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder19_zero	:	STD_LOGIC;
	 COMPONENT  prueba1_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder19_w_lg_zero1318w & wire_altpriority_encoder19_w_lg_w_lg_zero1320w1321w);
	zero <= (wire_altpriority_encoder18_zero AND wire_altpriority_encoder19_zero);
	altpriority_encoder18 :  prueba1_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder18_q,
		zero => wire_altpriority_encoder18_zero
	  );
	loop120 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder19_w_lg_w_lg_zero1318w1319w(i) <= wire_altpriority_encoder19_w_lg_zero1318w(0) AND wire_altpriority_encoder19_q(i);
	END GENERATE loop120;
	loop121 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder19_w_lg_zero1320w(i) <= wire_altpriority_encoder19_zero AND wire_altpriority_encoder18_q(i);
	END GENERATE loop121;
	wire_altpriority_encoder19_w_lg_zero1318w(0) <= NOT wire_altpriority_encoder19_zero;
	loop122 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder19_w_lg_w_lg_zero1320w1321w(i) <= wire_altpriority_encoder19_w_lg_zero1320w(i) OR wire_altpriority_encoder19_w_lg_w_lg_zero1318w1319w(i);
	END GENERATE loop122;
	altpriority_encoder19 :  prueba1_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder19_q,
		zero => wire_altpriority_encoder19_zero
	  );

 END RTL; --prueba1_altpriority_encoder_be8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altpriority_encoder_r08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END prueba1_altpriority_encoder_r08;

 ARCHITECTURE RTL OF prueba1_altpriority_encoder_r08 IS

	 SIGNAL  wire_altpriority_encoder10_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_w_lg_zero1272w1273w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_zero1274w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_zero1272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_w_lg_w_lg_zero1274w1275w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_zero	:	STD_LOGIC;
	 COMPONENT  prueba1_altpriority_encoder_bv7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder11_w_lg_zero1272w & wire_altpriority_encoder11_w_lg_w_lg_zero1274w1275w);
	altpriority_encoder10 :  prueba1_altpriority_encoder_bv7
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder10_q
	  );
	loop123 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder11_w_lg_w_lg_zero1272w1273w(i) <= wire_altpriority_encoder11_w_lg_zero1272w(0) AND wire_altpriority_encoder11_q(i);
	END GENERATE loop123;
	loop124 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder11_w_lg_zero1274w(i) <= wire_altpriority_encoder11_zero AND wire_altpriority_encoder10_q(i);
	END GENERATE loop124;
	wire_altpriority_encoder11_w_lg_zero1272w(0) <= NOT wire_altpriority_encoder11_zero;
	loop125 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder11_w_lg_w_lg_zero1274w1275w(i) <= wire_altpriority_encoder11_w_lg_zero1274w(i) OR wire_altpriority_encoder11_w_lg_w_lg_zero1272w1273w(i);
	END GENERATE loop125;
	altpriority_encoder11 :  prueba1_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder11_q,
		zero => wire_altpriority_encoder11_zero
	  );

 END RTL; --prueba1_altpriority_encoder_r08


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q zero
--VERSION_BEGIN 15.1 cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altpriority_encoder_rf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END prueba1_altpriority_encoder_rf8;

 ARCHITECTURE RTL OF prueba1_altpriority_encoder_rf8 IS

	 SIGNAL  wire_altpriority_encoder20_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder21_w_lg_w_lg_zero1328w1329w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_w_lg_zero1330w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_w_lg_zero1328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_w_lg_w_lg_zero1330w1331w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_zero	:	STD_LOGIC;
	 COMPONENT  prueba1_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder21_w_lg_zero1328w & wire_altpriority_encoder21_w_lg_w_lg_zero1330w1331w);
	zero <= (wire_altpriority_encoder20_zero AND wire_altpriority_encoder21_zero);
	altpriority_encoder20 :  prueba1_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder20_q,
		zero => wire_altpriority_encoder20_zero
	  );
	loop126 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder21_w_lg_w_lg_zero1328w1329w(i) <= wire_altpriority_encoder21_w_lg_zero1328w(0) AND wire_altpriority_encoder21_q(i);
	END GENERATE loop126;
	loop127 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder21_w_lg_zero1330w(i) <= wire_altpriority_encoder21_zero AND wire_altpriority_encoder20_q(i);
	END GENERATE loop127;
	wire_altpriority_encoder21_w_lg_zero1328w(0) <= NOT wire_altpriority_encoder21_zero;
	loop128 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder21_w_lg_w_lg_zero1330w1331w(i) <= wire_altpriority_encoder21_w_lg_zero1330w(i) OR wire_altpriority_encoder21_w_lg_w_lg_zero1328w1329w(i);
	END GENERATE loop128;
	altpriority_encoder21 :  prueba1_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder21_q,
		zero => wire_altpriority_encoder21_zero
	  );

 END RTL; --prueba1_altpriority_encoder_rf8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altpriority_encoder_tv8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END prueba1_altpriority_encoder_tv8;

 ARCHITECTURE RTL OF prueba1_altpriority_encoder_tv8 IS

	 SIGNAL  wire_altpriority_encoder8_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_w_lg_zero1263w1264w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_zero1265w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_zero1263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_w_lg_w_lg_zero1265w1266w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder9_zero	:	STD_LOGIC;
	 COMPONENT  prueba1_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder9_w_lg_zero1263w & wire_altpriority_encoder9_w_lg_w_lg_zero1265w1266w);
	altpriority_encoder8 :  prueba1_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder8_q
	  );
	loop129 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder9_w_lg_w_lg_zero1263w1264w(i) <= wire_altpriority_encoder9_w_lg_zero1263w(0) AND wire_altpriority_encoder9_q(i);
	END GENERATE loop129;
	loop130 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder9_w_lg_zero1265w(i) <= wire_altpriority_encoder9_zero AND wire_altpriority_encoder8_q(i);
	END GENERATE loop130;
	wire_altpriority_encoder9_w_lg_zero1263w(0) <= NOT wire_altpriority_encoder9_zero;
	loop131 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder9_w_lg_w_lg_zero1265w1266w(i) <= wire_altpriority_encoder9_w_lg_zero1265w(i) OR wire_altpriority_encoder9_w_lg_w_lg_zero1263w1264w(i);
	END GENERATE loop131;
	altpriority_encoder9 :  prueba1_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder9_q,
		zero => wire_altpriority_encoder9_zero
	  );

 END RTL; --prueba1_altpriority_encoder_tv8


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" PIPELINE=0 WIDTH=32 WIDTHAD=5 data q zero
--VERSION_BEGIN 15.1 cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altpriority_encoder_te9 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END prueba1_altpriority_encoder_te9;

 ARCHITECTURE RTL OF prueba1_altpriority_encoder_te9 IS

	 SIGNAL  wire_altpriority_encoder22_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder23_w_lg_w_lg_zero1338w1339w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_w_lg_zero1340w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_w_lg_zero1338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_w_lg_w_lg_zero1340w1341w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder23_zero	:	STD_LOGIC;
	 COMPONENT  prueba1_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder23_w_lg_zero1338w & wire_altpriority_encoder23_w_lg_w_lg_zero1340w1341w);
	zero <= (wire_altpriority_encoder22_zero AND wire_altpriority_encoder23_zero);
	altpriority_encoder22 :  prueba1_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder22_q,
		zero => wire_altpriority_encoder22_zero
	  );
	loop132 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder23_w_lg_w_lg_zero1338w1339w(i) <= wire_altpriority_encoder23_w_lg_zero1338w(0) AND wire_altpriority_encoder23_q(i);
	END GENERATE loop132;
	loop133 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder23_w_lg_zero1340w(i) <= wire_altpriority_encoder23_zero AND wire_altpriority_encoder22_q(i);
	END GENERATE loop133;
	wire_altpriority_encoder23_w_lg_zero1338w(0) <= NOT wire_altpriority_encoder23_zero;
	loop134 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder23_w_lg_w_lg_zero1340w1341w(i) <= wire_altpriority_encoder23_w_lg_zero1340w(i) OR wire_altpriority_encoder23_w_lg_w_lg_zero1338w1339w(i);
	END GENERATE loop134;
	altpriority_encoder23 :  prueba1_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder23_q,
		zero => wire_altpriority_encoder23_zero
	  );

 END RTL; --prueba1_altpriority_encoder_te9

--synthesis_resources = reg 6 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altpriority_encoder_uja IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0)
	 ); 
 END prueba1_altpriority_encoder_uja;

 ARCHITECTURE RTL OF prueba1_altpriority_encoder_uja IS

	 SIGNAL  wire_altpriority_encoder6_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_w_lg_zero1253w1254w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_zero1255w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_zero1253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_w_lg_w_lg_zero1255w1256w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder7_zero	:	STD_LOGIC;
	 SIGNAL	 pipeline_q_dffe	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  tmp_q_wire :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 COMPONENT  prueba1_altpriority_encoder_tv8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altpriority_encoder_te9
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= pipeline_q_dffe;
	tmp_q_wire <= ( wire_altpriority_encoder7_w_lg_zero1253w & wire_altpriority_encoder7_w_lg_w_lg_zero1255w1256w);
	altpriority_encoder6 :  prueba1_altpriority_encoder_tv8
	  PORT MAP ( 
		data => data(31 DOWNTO 0),
		q => wire_altpriority_encoder6_q
	  );
	loop135 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder7_w_lg_w_lg_zero1253w1254w(i) <= wire_altpriority_encoder7_w_lg_zero1253w(0) AND wire_altpriority_encoder7_q(i);
	END GENERATE loop135;
	loop136 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder7_w_lg_zero1255w(i) <= wire_altpriority_encoder7_zero AND wire_altpriority_encoder6_q(i);
	END GENERATE loop136;
	wire_altpriority_encoder7_w_lg_zero1253w(0) <= NOT wire_altpriority_encoder7_zero;
	loop137 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder7_w_lg_w_lg_zero1255w1256w(i) <= wire_altpriority_encoder7_w_lg_zero1255w(i) OR wire_altpriority_encoder7_w_lg_w_lg_zero1253w1254w(i);
	END GENERATE loop137;
	altpriority_encoder7 :  prueba1_altpriority_encoder_te9
	  PORT MAP ( 
		data => data(63 DOWNTO 32),
		q => wire_altpriority_encoder7_q,
		zero => wire_altpriority_encoder7_zero
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN pipeline_q_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN pipeline_q_dffe <= tmp_q_wire;
			END IF;
		END IF;
	END PROCESS;

 END RTL; --prueba1_altpriority_encoder_uja


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 15.1 cbx_altpriority_encoder 2015:10:21:18:09:23:SJ cbx_mgl 2015:10:21:18:12:49:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altpriority_encoder_q08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END prueba1_altpriority_encoder_q08;

 ARCHITECTURE RTL OF prueba1_altpriority_encoder_q08 IS

	 SIGNAL  wire_altpriority_encoder24_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_w_lg_w_lg_zero1348w1349w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_w_lg_zero1350w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_w_lg_zero1348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_w_lg_w_lg_zero1350w1351w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder25_zero	:	STD_LOGIC;
	 COMPONENT  prueba1_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder25_w_lg_zero1348w & wire_altpriority_encoder25_w_lg_w_lg_zero1350w1351w);
	altpriority_encoder24 :  prueba1_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder24_q
	  );
	loop138 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder25_w_lg_w_lg_zero1348w1349w(i) <= wire_altpriority_encoder25_w_lg_zero1348w(0) AND wire_altpriority_encoder25_q(i);
	END GENERATE loop138;
	loop139 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder25_w_lg_zero1350w(i) <= wire_altpriority_encoder25_zero AND wire_altpriority_encoder24_q(i);
	END GENERATE loop139;
	wire_altpriority_encoder25_w_lg_zero1348w(0) <= NOT wire_altpriority_encoder25_zero;
	loop140 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder25_w_lg_w_lg_zero1350w1351w(i) <= wire_altpriority_encoder25_w_lg_zero1350w(i) OR wire_altpriority_encoder25_w_lg_w_lg_zero1348w1349w(i);
	END GENERATE loop140;
	altpriority_encoder25 :  prueba1_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder25_q,
		zero => wire_altpriority_encoder25_zero
	  );

 END RTL; --prueba1_altpriority_encoder_q08

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = altsquare 1 lpm_add_sub 42 lpm_mult 5 lpm_mux 5 mux21 31 reg 1569 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  prueba1_altfp_log_8ka IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END prueba1_altfp_log_8ka;

 ARCHITECTURE RTL OF prueba1_altfp_log_8ka IS

	 SIGNAL  wire_Lshiftsmall_data	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Lshiftsmall_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_data	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_distance	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_E_w_lg_q189w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_L_result	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_data	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_Rshiftsmall_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_exp_nan_result	:	STD_LOGIC;
	 SIGNAL  wire_exp_zero_result	:	STD_LOGIC;
	 SIGNAL  wire_man_inf_result	:	STD_LOGIC;
	 SIGNAL  wire_man_nan_result	:	STD_LOGIC;
	 SIGNAL  wire_add1_dataa	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add1_result	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add2_dataa	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add2_datab	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add2_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_exp_biase_sub_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_sub1_dataa	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_sub1_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_sub2_dataa	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_sub2_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_sub3_dataa	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_sub3_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_sub3_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_sub4_datab	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_sub4_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_sub5_dataa	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_sub5_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_sub5_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_sub6_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_sub6_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_range_reduction_almostlog	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_range_reduction_z	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_E_data	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_lzc_norm_E_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_lzoc_data	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_lzoc_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_squarer_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL	 absELog2_pipe_reg0	:	STD_LOGIC_VECTOR(34 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absELog2_pipe_reg1	:	STD_LOGIC_VECTOR(34 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absELog2_pipe_reg2	:	STD_LOGIC_VECTOR(34 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg0	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg1	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg2	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg3	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg4	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg5	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg6	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg7	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg8	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0_pipe_reg9	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0s_pipe1_reg0	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0s_pipe1_reg1	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0s_pipe1_reg2	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0s_pipe1_reg3	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 absZ0s_reg0	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 almostLog_pipe_reg0	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 almostLog_pipe_reg1	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 almostLog_pipe_reg2	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 doRR_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 doRR_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg0	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg1	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg2	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg3	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg4	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg5	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg6	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg7	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg8	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E0_pipe_reg9	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 E_normal_pipe_reg0	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_is_ebiase_pipe_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_is_ebiase_pipe_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_is_ebiase_pipe_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg10	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg11	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg12	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg13	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg14	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg15	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg16	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg17	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg5	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg6	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg7	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg8	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_infinity_pipe_reg9	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg10	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg11	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg12	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg13	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg14	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg15	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg16	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg17	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg5	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg6	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg7	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg8	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_nan_pipe_reg9	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg10	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg11	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg12	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg13	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg14	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg15	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg16	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg17	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg5	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg6	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg7	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg8	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_one_pipe_reg9	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg10	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg11	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg12	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg13	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg14	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg15	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg16	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg17	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg5	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg6	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg7	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg8	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_is_zero_pipe_reg9	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Log_normal_normd_pipe_reg0	:	STD_LOGIC_VECTOR(46 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Log_normal_reg0	:	STD_LOGIC_VECTOR(46 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Log_small_normd_pipe_reg0	:	STD_LOGIC_VECTOR(26 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Log_small_normd_pipe_reg1	:	STD_LOGIC_VECTOR(26 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Lshiftval_reg0	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Lshiftval_reg1	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Lshiftval_reg2	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Lshiftval_reg3	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg0	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg1	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg2	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg3	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg4	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg5	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg6	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg7	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg8	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_pipe1_reg9	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg0	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg1	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg2	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg3	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg4	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg5	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg6	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 lzo_reg7	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_data_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_data_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_data_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg5	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg6	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg7	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg8	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 small_flag_pipe_reg9	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg5	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg6	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg7	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg8	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe1_reg9	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe2_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe2_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe2_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe2_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe2_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe2_reg5	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe3_reg0	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe3_reg1	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe3_reg2	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe3_reg3	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sR_pipe3_reg4	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Z2o2_pipe_reg0	:	STD_LOGIC_VECTOR(13 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Z2o2_small_s_pipe_reg0	:	STD_LOGIC_VECTOR(13 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Zfinal_reg0	:	STD_LOGIC_VECTOR(25 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Zfinal_reg1	:	STD_LOGIC_VECTOR(25 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_addsub1_result	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_addsub2_add_sub	:	STD_LOGIC;
	 SIGNAL  wire_addsub2_result	:	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  wire_mult1_result	:	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL	wire_mux_result0a_dataout	:	STD_LOGIC_VECTOR(30 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_doRR_pipe125w126w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_First_bit9w83w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_small_flag206w215w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_small_flag206w207w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sR_pipe188w89w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sR_pipe292w93w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_E0_range42w43w44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_E0_range46w47w48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_E0_range50w51w52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_E0_range54w55w56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_E0_range58w59w60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_E0_range62w63w64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_E0_range66w67w68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_exp_data_range31w33w34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_Log_small_range149w154w194w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_Log_small_range150w198w199w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_sR254w255w256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_doRR_pipe124w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_w_lg_First_bit82w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_w_lg_small_flag214w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_small_flag204w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_lg_sR_pipe187w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_w_lg_sR_pipe291w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_range13w15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_range16w18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_range19w21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_range22w24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_range25w27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_range28w30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_g_range228w229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_small_range149w192w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_small_range150w197w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_lg_doRR111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_doRR_pipe125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_E_normal212w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_all_zero240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_First_bit9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_is_one247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_man_all_zero241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_small_flag206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sR_pipe188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sR_pipe292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sR_pipe3179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range38w39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range42w43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range46w47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range50w51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range54w55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range58w59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range62w63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_E0_range66w67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_data_range31w33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_small_range149w154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_small_range150w198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_input_is_one247w248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_input_is_zero244w245w246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_input_is_zero244w245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_sR254w255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_input_is_zero244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sR254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_g_range220w221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_g_range223w224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_g_range226w227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_small_range150w155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_Log_small_range150w151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_First_bit96w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  absE :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  absELog2 :	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  absELog2_pad :	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  absELog2_pipe :	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  absZ0 :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  absZ0_pipe :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  absZ0s :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  absZ0s_pipe1 :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  absZ0s_pipe2 :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  almostLog :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  almostLog_pipe :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  data_exp_is_ebiase :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  doRR :	STD_LOGIC;
	 SIGNAL  doRR_pipe :	STD_LOGIC;
	 SIGNAL  E0 :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  E0_is_zero :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  E0_pipe :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  E0_sub :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  E0offset :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  E_normal :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  E_normal_pipe :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  E_small :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  EFR :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  ER :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_all_one :	STD_LOGIC;
	 SIGNAL  exp_all_zero :	STD_LOGIC;
	 SIGNAL  exp_biase :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_data :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_is_ebiase :	STD_LOGIC;
	 SIGNAL  exp_is_ebiase_pipe :	STD_LOGIC;
	 SIGNAL  First_bit :	STD_LOGIC;
	 SIGNAL  input_is_infinity :	STD_LOGIC;
	 SIGNAL  input_is_infinity_pipe :	STD_LOGIC;
	 SIGNAL  input_is_nan :	STD_LOGIC;
	 SIGNAL  input_is_nan_pipe :	STD_LOGIC;
	 SIGNAL  input_is_one :	STD_LOGIC;
	 SIGNAL  input_is_one_pipe :	STD_LOGIC;
	 SIGNAL  input_is_zero :	STD_LOGIC;
	 SIGNAL  input_is_zero_pipe :	STD_LOGIC;
	 SIGNAL  Log1p_normal :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  Log2 :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Log_g :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Log_normal :	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  Log_normal_normd :	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  Log_normal_normd_pipe :	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  Log_normal_pipe :	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  Log_small :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  Log_small1 :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Log_small2 :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Log_small_normd :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Log_small_normd_pipe :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  LogF_normal :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  LogF_normal_pad :	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  Lshiftval :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  lzo :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  lzo_pipe1 :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  lzo_pipe2 :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  man_above_half :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  man_all_zero :	STD_LOGIC;
	 SIGNAL  man_below_half :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  man_data :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_not_zero :	STD_LOGIC;
	 SIGNAL  pfinal_s :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  round :	STD_LOGIC;
	 SIGNAL  Rshiftval :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  sign_data :	STD_LOGIC;
	 SIGNAL  sign_data_pipe :	STD_LOGIC;
	 SIGNAL  small_flag :	STD_LOGIC;
	 SIGNAL  small_flag_pipe :	STD_LOGIC;
	 SIGNAL  squarerIn :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  squarerIn0 :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  squarerIn1 :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  sR :	STD_LOGIC;
	 SIGNAL  sR_pipe1 :	STD_LOGIC;
	 SIGNAL  sR_pipe2 :	STD_LOGIC;
	 SIGNAL  sR_pipe3 :	STD_LOGIC;
	 SIGNAL  sticky :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w203w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Y0 :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Z2o2 :	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  Z2o2_pipe :	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  Z2o2_small :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  Z2o2_small_s :	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  Z2o2_small_s_pipe :	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  Z_small :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  Zfinal :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  Zfinal_pipe :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_w_data_exp_is_ebiase_range6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_exp_is_ebiase_range14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_exp_is_ebiase_range17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_exp_is_ebiase_range20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_exp_is_ebiase_range23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_exp_is_ebiase_range26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_exp_is_ebiase_range29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_range66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_is_zero_range40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_is_zero_range45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_is_zero_range49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_is_zero_range53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_is_zero_range57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_is_zero_range61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_E0_is_zero_range65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_range13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_range16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_range19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_range22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_range25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_range28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_data_range31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_Log_g_range220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_Log_g_range223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_Log_g_range228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_Log_g_range226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_Log_normal_normd_range205w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_Log_small_range193w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_Log_small_range191w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_Log_small_range149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_Log_small_range196w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_w_Log_small_range150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_range218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_range222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_range225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_Y0_range86w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_w_Y0_range95w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 COMPONENT  prueba1_altbarrel_shift_05e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altbarrel_shift_8ib
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(5 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(63 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altbarrel_shift_j8e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		distance	:	IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		result	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_and_or_f9b
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_and_or_t6b
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_and_or_a8b
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(22 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_csa_s0e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(38 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(38 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(38 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_csa_k0e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(30 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(30 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(30 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_csa_0nc
	 PORT
	 ( 
		dataa	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_csa_d4b
	 PORT
	 ( 
		dataa	:	IN  STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(11 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_csa_umc
	 PORT
	 ( 
		dataa	:	IN  STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_csa_nlf
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(25 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(25 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altfp_log_csa_8kf
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(7 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_range_reduction_c2e
	 PORT
	 ( 
		a0_in	:	IN  STD_LOGIC_VECTOR(4 DOWNTO 0);
		aclr	:	IN  STD_LOGIC := '0';
		almostlog	:	OUT  STD_LOGIC_VECTOR(38 DOWNTO 0);
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC;
		y0_in	:	IN  STD_LOGIC_VECTOR(24 DOWNTO 0);
		z	:	OUT  STD_LOGIC_VECTOR(25 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altpriority_encoder_uja
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clk_en	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  prueba1_altpriority_encoder_q08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  altsquare
	 GENERIC 
	 (
		DATA_WIDTH	:	NATURAL;
		PIPELINE	:	NATURAL;
		REPRESENTATION	:	STRING := "UNSIGNED";
		RESULT_ALIGNMENT	:	STRING := "LSB";
		RESULT_WIDTH	:	NATURAL;
		lpm_type	:	STRING := "altsquare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clock	:	IN STD_LOGIC := '1';
		data	:	IN STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
		ena	:	IN STD_LOGIC := '1';
		result	:	OUT STD_LOGIC_VECTOR(RESULT_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop141 : FOR i IN 0 TO 12 GENERATE 
		wire_w_lg_w_lg_doRR_pipe125w126w(i) <= wire_w_lg_doRR_pipe125w(0) AND squarerIn0(i);
	END GENERATE loop141;
	loop142 : FOR i IN 0 TO 24 GENERATE 
		wire_w_lg_w_lg_First_bit9w83w(i) <= wire_w_lg_First_bit9w(0) AND man_below_half(i);
	END GENERATE loop142;
	loop143 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_small_flag206w215w(i) <= wire_w_lg_small_flag206w(0) AND wire_sub6_result(i);
	END GENERATE loop143;
	loop144 : FOR i IN 0 TO 26 GENERATE 
		wire_w_lg_w_lg_small_flag206w207w(i) <= wire_w_lg_small_flag206w(0) AND wire_w_Log_normal_normd_range205w(i);
	END GENERATE loop144;
	loop145 : FOR i IN 0 TO 11 GENERATE 
		wire_w_lg_w_lg_sR_pipe188w89w(i) <= wire_w_lg_sR_pipe188w(0) AND wire_w_Y0_range86w(i);
	END GENERATE loop145;
	loop146 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_sR_pipe292w93w(i) <= wire_w_lg_sR_pipe292w(0) AND E0(i);
	END GENERATE loop146;
	wire_w_lg_w_lg_w_E0_range42w43w44w(0) <= wire_w_lg_w_E0_range42w43w(0) AND wire_w_E0_is_zero_range40w(0);
	wire_w_lg_w_lg_w_E0_range46w47w48w(0) <= wire_w_lg_w_E0_range46w47w(0) AND wire_w_E0_is_zero_range45w(0);
	wire_w_lg_w_lg_w_E0_range50w51w52w(0) <= wire_w_lg_w_E0_range50w51w(0) AND wire_w_E0_is_zero_range49w(0);
	wire_w_lg_w_lg_w_E0_range54w55w56w(0) <= wire_w_lg_w_E0_range54w55w(0) AND wire_w_E0_is_zero_range53w(0);
	wire_w_lg_w_lg_w_E0_range58w59w60w(0) <= wire_w_lg_w_E0_range58w59w(0) AND wire_w_E0_is_zero_range57w(0);
	wire_w_lg_w_lg_w_E0_range62w63w64w(0) <= wire_w_lg_w_E0_range62w63w(0) AND wire_w_E0_is_zero_range61w(0);
	wire_w_lg_w_lg_w_E0_range66w67w68w(0) <= wire_w_lg_w_E0_range66w67w(0) AND wire_w_E0_is_zero_range65w(0);
	wire_w_lg_w_lg_w_exp_data_range31w33w34w(0) <= wire_w_lg_w_exp_data_range31w33w(0) AND wire_w_data_exp_is_ebiase_range29w(0);
	loop147 : FOR i IN 0 TO 26 GENERATE 
		wire_w_lg_w_lg_w_Log_small_range149w154w194w(i) <= wire_w_lg_w_Log_small_range149w154w(0) AND wire_w_Log_small_range193w(i);
	END GENERATE loop147;
	loop148 : FOR i IN 0 TO 26 GENERATE 
		wire_w_lg_w_lg_w_Log_small_range150w198w199w(i) <= wire_w_lg_w_Log_small_range150w198w(0) AND Log_small1(i);
	END GENERATE loop148;
	wire_w_lg_w_lg_w_lg_sR254w255w256w(0) <= wire_w_lg_w_lg_sR254w255w(0) AND wire_w_lg_input_is_one247w(0);
	loop149 : FOR i IN 0 TO 12 GENERATE 
		wire_w_lg_doRR_pipe124w(i) <= doRR_pipe AND squarerIn1(i);
	END GENERATE loop149;
	loop150 : FOR i IN 0 TO 24 GENERATE 
		wire_w_lg_First_bit82w(i) <= First_bit AND man_above_half(i);
	END GENERATE loop150;
	loop151 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_small_flag214w(i) <= small_flag AND E_small(i);
	END GENERATE loop151;
	loop152 : FOR i IN 0 TO 26 GENERATE 
		wire_w_lg_small_flag204w(i) <= small_flag AND wire_w203w(i);
	END GENERATE loop152;
	loop153 : FOR i IN 0 TO 11 GENERATE 
		wire_w_lg_sR_pipe187w(i) <= sR_pipe1 AND wire_sub1_result(i);
	END GENERATE loop153;
	loop154 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_sR_pipe291w(i) <= sR_pipe2 AND wire_sub2_result(i);
	END GENERATE loop154;
	wire_w_lg_w_exp_data_range13w15w(0) <= wire_w_exp_data_range13w(0) AND wire_w_data_exp_is_ebiase_range6w(0);
	wire_w_lg_w_exp_data_range16w18w(0) <= wire_w_exp_data_range16w(0) AND wire_w_data_exp_is_ebiase_range14w(0);
	wire_w_lg_w_exp_data_range19w21w(0) <= wire_w_exp_data_range19w(0) AND wire_w_data_exp_is_ebiase_range17w(0);
	wire_w_lg_w_exp_data_range22w24w(0) <= wire_w_exp_data_range22w(0) AND wire_w_data_exp_is_ebiase_range20w(0);
	wire_w_lg_w_exp_data_range25w27w(0) <= wire_w_exp_data_range25w(0) AND wire_w_data_exp_is_ebiase_range23w(0);
	wire_w_lg_w_exp_data_range28w30w(0) <= wire_w_exp_data_range28w(0) AND wire_w_data_exp_is_ebiase_range26w(0);
	wire_w_lg_w_Log_g_range228w229w(0) <= wire_w_Log_g_range228w(0) AND wire_w_lg_w_Log_g_range226w227w(0);
	loop155 : FOR i IN 0 TO 26 GENERATE 
		wire_w_lg_w_Log_small_range149w192w(i) <= wire_w_Log_small_range149w(0) AND wire_w_Log_small_range191w(i);
	END GENERATE loop155;
	loop156 : FOR i IN 0 TO 26 GENERATE 
		wire_w_lg_w_Log_small_range150w197w(i) <= wire_w_Log_small_range150w(0) AND wire_w_Log_small_range196w(i);
	END GENERATE loop156;
	wire_w_lg_doRR111w(0) <= NOT doRR;
	wire_w_lg_doRR_pipe125w(0) <= NOT doRR_pipe;
	loop157 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_E_normal212w(i) <= NOT E_normal(i);
	END GENERATE loop157;
	wire_w_lg_exp_all_zero240w(0) <= NOT exp_all_zero;
	wire_w_lg_First_bit9w(0) <= NOT First_bit;
	wire_w_lg_input_is_one247w(0) <= NOT input_is_one;
	wire_w_lg_man_all_zero241w(0) <= NOT man_all_zero;
	wire_w_lg_small_flag206w(0) <= NOT small_flag;
	wire_w_lg_sR_pipe188w(0) <= NOT sR_pipe1;
	wire_w_lg_sR_pipe292w(0) <= NOT sR_pipe2;
	wire_w_lg_sR_pipe3179w(0) <= NOT sR_pipe3;
	wire_w_lg_w_E0_range38w39w(0) <= NOT wire_w_E0_range38w(0);
	wire_w_lg_w_E0_range42w43w(0) <= NOT wire_w_E0_range42w(0);
	wire_w_lg_w_E0_range46w47w(0) <= NOT wire_w_E0_range46w(0);
	wire_w_lg_w_E0_range50w51w(0) <= NOT wire_w_E0_range50w(0);
	wire_w_lg_w_E0_range54w55w(0) <= NOT wire_w_E0_range54w(0);
	wire_w_lg_w_E0_range58w59w(0) <= NOT wire_w_E0_range58w(0);
	wire_w_lg_w_E0_range62w63w(0) <= NOT wire_w_E0_range62w(0);
	wire_w_lg_w_E0_range66w67w(0) <= NOT wire_w_E0_range66w(0);
	wire_w_lg_w_exp_data_range31w33w(0) <= NOT wire_w_exp_data_range31w(0);
	wire_w_lg_w_Log_small_range149w154w(0) <= NOT wire_w_Log_small_range149w(0);
	wire_w_lg_w_Log_small_range150w198w(0) <= NOT wire_w_Log_small_range150w(0);
	wire_w_lg_w_lg_input_is_one247w248w(0) <= wire_w_lg_input_is_one247w(0) OR input_is_nan;
	wire_w_lg_w_lg_w_lg_input_is_zero244w245w246w(0) <= wire_w_lg_w_lg_input_is_zero244w245w(0) OR input_is_one;
	wire_w_lg_w_lg_input_is_zero244w245w(0) <= wire_w_lg_input_is_zero244w(0) OR input_is_nan;
	wire_w_lg_w_lg_sR254w255w(0) <= wire_w_lg_sR254w(0) OR input_is_nan;
	wire_w_lg_input_is_zero244w(0) <= input_is_zero OR input_is_infinity;
	wire_w_lg_sR254w(0) <= sR OR input_is_zero;
	wire_w_lg_w_Log_g_range220w221w(0) <= wire_w_Log_g_range220w(0) OR wire_w_sticky_range218w(0);
	wire_w_lg_w_Log_g_range223w224w(0) <= wire_w_Log_g_range223w(0) OR wire_w_sticky_range222w(0);
	wire_w_lg_w_Log_g_range226w227w(0) <= wire_w_Log_g_range226w(0) OR wire_w_sticky_range225w(0);
	wire_w_lg_w_Log_small_range150w155w(0) <= wire_w_Log_small_range150w(0) OR wire_w_lg_w_Log_small_range149w154w(0);
	wire_w_lg_w_Log_small_range150w151w(0) <= wire_w_Log_small_range150w(0) OR wire_w_Log_small_range149w(0);
	loop158 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_First_bit96w(i) <= First_bit XOR wire_w_Y0_range95w(i);
	END GENERATE loop158;
	absE <= (wire_w_lg_w_lg_sR_pipe292w93w OR wire_w_lg_sR_pipe291w);
	absELog2 <= absELog2_pipe_reg2;
	absELog2_pad <= ( absELog2 & "000000000000");
	absELog2_pipe <= wire_mult1_result;
	absZ0 <= absZ0_pipe_reg9;
	absZ0_pipe <= (wire_w_lg_w_lg_sR_pipe188w89w OR wire_w_lg_sR_pipe187w);
	absZ0s <= wire_Lshiftsmall_result(31 DOWNTO 20);
	absZ0s_pipe1 <= absZ0s_reg0;
	absZ0s_pipe2 <= absZ0s_pipe1_reg3;
	aclr <= '0';
	almostLog <= almostLog_pipe_reg2;
	almostLog_pipe <= wire_range_reduction_almostlog;
	clk_en <= '1';
	data_exp_is_ebiase <= ( wire_w_lg_w_lg_w_exp_data_range31w33w34w & wire_w_lg_w_exp_data_range28w30w & wire_w_lg_w_exp_data_range25w27w & wire_w_lg_w_exp_data_range22w24w & wire_w_lg_w_exp_data_range19w21w & wire_w_lg_w_exp_data_range16w18w & wire_w_lg_w_exp_data_range13w15w & exp_data(0));
	doRR <= Lshiftval(5);
	doRR_pipe <= doRR_reg1(0);
	E0 <= E0_pipe_reg9;
	E0_is_zero <= ( wire_w_lg_w_lg_w_E0_range66w67w68w & wire_w_lg_w_lg_w_E0_range62w63w64w & wire_w_lg_w_lg_w_E0_range58w59w60w & wire_w_lg_w_lg_w_E0_range54w55w56w & wire_w_lg_w_lg_w_E0_range50w51w52w & wire_w_lg_w_lg_w_E0_range46w47w48w & wire_w_lg_w_lg_w_E0_range42w43w44w & wire_w_lg_w_E0_range38w39w);
	E0_pipe <= wire_exp_biase_sub_result;
	E0_sub <= ( wire_w_lg_w_Log_small_range150w151w & wire_w_lg_w_Log_small_range150w155w);
	E0offset <= "10000110";
	E_normal <= E_normal_pipe_reg0;
	E_normal_pipe <= wire_lzc_norm_E_q(4 DOWNTO 0);
	E_small <= wire_sub5_result;
	EFR <= wire_add2_result;
	ER <= (wire_w_lg_w_lg_small_flag206w215w OR wire_w_lg_small_flag214w);
	exp_all_one <= wire_exp_nan_result;
	exp_all_zero <= wire_exp_zero_result;
	exp_biase <= ( "0111111" & wire_w_lg_First_bit9w);
	exp_data <= data(30 DOWNTO 23);
	exp_is_ebiase <= exp_is_ebiase_pipe_reg2(0);
	exp_is_ebiase_pipe <= data_exp_is_ebiase(7);
	First_bit <= man_data(22);
	input_is_infinity <= input_is_infinity_pipe_reg17(0);
	input_is_infinity_pipe <= (exp_all_one AND wire_w_lg_man_all_zero241w(0));
	input_is_nan <= input_is_nan_pipe_reg17(0);
	input_is_nan_pipe <= ((exp_all_one AND man_not_zero) OR sign_data_pipe);
	input_is_one <= input_is_one_pipe_reg17(0);
	input_is_one_pipe <= (exp_is_ebiase AND wire_w_lg_man_all_zero241w(0));
	input_is_zero <= input_is_zero_pipe_reg17(0);
	input_is_zero_pipe <= wire_w_lg_exp_all_zero240w(0);
	Log1p_normal <= wire_sub4_result;
	Log2 <= "101100010111001000011000000";
	Log_g <= (wire_w_lg_w_lg_small_flag206w207w OR wire_w_lg_small_flag204w);
	Log_normal <= wire_addsub2_result;
	Log_normal_normd <= Log_normal_normd_pipe_reg0;
	Log_normal_normd_pipe <= wire_lzc_norm_L_result(63 DOWNTO 17);
	Log_normal_pipe <= Log_normal_reg0;
	Log_small <= wire_addsub1_result;
	Log_small1 <= (wire_w_lg_w_lg_w_Log_small_range149w154w194w OR wire_w_lg_w_Log_small_range149w192w);
	Log_small2 <= (wire_w_lg_w_lg_w_Log_small_range150w198w199w OR wire_w_lg_w_Log_small_range150w197w);
	Log_small_normd <= Log_small_normd_pipe_reg1;
	Log_small_normd_pipe <= Log_small2;
	LogF_normal <= wire_add1_result;
	LogF_normal_pad <= ( LogF_normal(38) & LogF_normal(38) & LogF_normal(38) & LogF_normal(38) & LogF_normal(38) & LogF_normal(38) & LogF_normal(38) & LogF_normal(38) & LogF_normal);
	Lshiftval <= wire_sub3_result;
	lzo <= lzo_pipe1_reg9;
	lzo_pipe1 <= (NOT wire_lzoc_q);
	lzo_pipe2 <= lzo_reg7;
	man_above_half <= ( "0" & "1" & man_data);
	man_all_zero <= wire_man_inf_result;
	man_below_half <= ( "1" & man_data & "0");
	man_data <= data(22 DOWNTO 0);
	man_not_zero <= wire_man_nan_result;
	pfinal_s <= "01101";
	result <= ( wire_w_lg_w_lg_w_lg_sR254w255w256w & wire_mux_result0a_dataout);
	round <= wire_w_lg_w_Log_g_range228w229w(0);
	Rshiftval <= Lshiftval_reg3;
	sign_data <= data(31);
	sign_data_pipe <= sign_data_reg2(0);
	small_flag <= small_flag_pipe_reg9(0);
	small_flag_pipe <= (wire_w_lg_doRR111w(0) AND E0_is_zero(7));
	squarerIn <= (wire_w_lg_w_lg_doRR_pipe125w126w OR wire_w_lg_doRR_pipe124w);
	squarerIn0 <= ( absZ0s_pipe1 & "0");
	squarerIn1 <= Zfinal(25 DOWNTO 13);
	sR <= sR_pipe3_reg4(0);
	sR_pipe1 <= (NOT (data_exp_is_ebiase(7) OR exp_data(7)));
	sR_pipe2 <= sR_pipe1_reg9(0);
	sR_pipe3 <= sR_pipe2_reg5(0);
	sticky <= ( wire_w_lg_w_Log_g_range223w224w & wire_w_lg_w_Log_g_range220w221w & Log_g(0));
	wire_w203w <= ( Log_small_normd(25 DOWNTO 0) & "0");
	Y0 <= (wire_w_lg_w_lg_First_bit9w83w OR wire_w_lg_First_bit82w);
	Z2o2 <= Z2o2_pipe_reg0;
	Z2o2_pipe <= wire_squarer_result;
	Z2o2_small <= ( "0000000000000" & Z2o2_small_s & "00");
	Z2o2_small_s <= Z2o2_small_s_pipe_reg0;
	Z2o2_small_s_pipe <= wire_Rshiftsmall_result(31 DOWNTO 18);
	Z_small <= ( absZ0s_pipe2 & "00000000000000000");
	Zfinal <= wire_range_reduction_z;
	Zfinal_pipe <= Zfinal_reg1;
	wire_w_data_exp_is_ebiase_range6w(0) <= data_exp_is_ebiase(0);
	wire_w_data_exp_is_ebiase_range14w(0) <= data_exp_is_ebiase(1);
	wire_w_data_exp_is_ebiase_range17w(0) <= data_exp_is_ebiase(2);
	wire_w_data_exp_is_ebiase_range20w(0) <= data_exp_is_ebiase(3);
	wire_w_data_exp_is_ebiase_range23w(0) <= data_exp_is_ebiase(4);
	wire_w_data_exp_is_ebiase_range26w(0) <= data_exp_is_ebiase(5);
	wire_w_data_exp_is_ebiase_range29w(0) <= data_exp_is_ebiase(6);
	wire_w_E0_range38w(0) <= E0(0);
	wire_w_E0_range42w(0) <= E0(1);
	wire_w_E0_range46w(0) <= E0(2);
	wire_w_E0_range50w(0) <= E0(3);
	wire_w_E0_range54w(0) <= E0(4);
	wire_w_E0_range58w(0) <= E0(5);
	wire_w_E0_range62w(0) <= E0(6);
	wire_w_E0_range66w(0) <= E0(7);
	wire_w_E0_is_zero_range40w(0) <= E0_is_zero(0);
	wire_w_E0_is_zero_range45w(0) <= E0_is_zero(1);
	wire_w_E0_is_zero_range49w(0) <= E0_is_zero(2);
	wire_w_E0_is_zero_range53w(0) <= E0_is_zero(3);
	wire_w_E0_is_zero_range57w(0) <= E0_is_zero(4);
	wire_w_E0_is_zero_range61w(0) <= E0_is_zero(5);
	wire_w_E0_is_zero_range65w(0) <= E0_is_zero(6);
	wire_w_exp_data_range13w(0) <= exp_data(1);
	wire_w_exp_data_range16w(0) <= exp_data(2);
	wire_w_exp_data_range19w(0) <= exp_data(3);
	wire_w_exp_data_range22w(0) <= exp_data(4);
	wire_w_exp_data_range25w(0) <= exp_data(5);
	wire_w_exp_data_range28w(0) <= exp_data(6);
	wire_w_exp_data_range31w(0) <= exp_data(7);
	wire_w_Log_g_range220w(0) <= Log_g(1);
	wire_w_Log_g_range223w(0) <= Log_g(2);
	wire_w_Log_g_range228w(0) <= Log_g(3);
	wire_w_Log_g_range226w(0) <= Log_g(4);
	wire_w_Log_normal_normd_range205w <= Log_normal_normd(45 DOWNTO 19);
	wire_w_Log_small_range193w <= Log_small(26 DOWNTO 0);
	wire_w_Log_small_range191w <= Log_small(27 DOWNTO 1);
	wire_w_Log_small_range149w(0) <= Log_small(27);
	wire_w_Log_small_range196w <= Log_small(28 DOWNTO 2);
	wire_w_Log_small_range150w(0) <= Log_small(28);
	wire_w_sticky_range218w(0) <= sticky(0);
	wire_w_sticky_range222w(0) <= sticky(1);
	wire_w_sticky_range225w(0) <= sticky(2);
	wire_w_Y0_range86w <= Y0(11 DOWNTO 0);
	wire_w_Y0_range95w <= Y0(23 DOWNTO 1);
	wire_Lshiftsmall_data <= ( absZ0 & "00000000000000000000");
	Lshiftsmall :  prueba1_altbarrel_shift_05e
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => wire_Lshiftsmall_data,
		distance => Lshiftval(4 DOWNTO 0),
		result => wire_Lshiftsmall_result
	  );
	wire_lzc_norm_L_data <= ( Log_normal_pipe & "00000000000000000");
	wire_lzc_norm_L_distance <= wire_lzc_norm_E_w_lg_q189w;
	loop159 : FOR i IN 0 TO 5 GENERATE 
		wire_lzc_norm_E_w_lg_q189w(i) <= NOT wire_lzc_norm_E_q(i);
	END GENERATE loop159;
	lzc_norm_L :  prueba1_altbarrel_shift_8ib
	  PORT MAP ( 
		data => wire_lzc_norm_L_data,
		distance => wire_lzc_norm_L_distance,
		result => wire_lzc_norm_L_result
	  );
	wire_Rshiftsmall_data <= ( Z2o2 & "000000000000000000");
	Rshiftsmall :  prueba1_altbarrel_shift_j8e
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => wire_Rshiftsmall_data,
		distance => Rshiftval(4 DOWNTO 0),
		result => wire_Rshiftsmall_result
	  );
	exp_nan :  prueba1_altfp_log_and_or_f9b
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => exp_data,
		result => wire_exp_nan_result
	  );
	exp_zero :  prueba1_altfp_log_and_or_t6b
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => exp_data,
		result => wire_exp_zero_result
	  );
	man_inf :  prueba1_altfp_log_and_or_a8b
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => man_data,
		result => wire_man_inf_result
	  );
	man_nan :  prueba1_altfp_log_and_or_a8b
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		data => man_data,
		result => wire_man_nan_result
	  );
	wire_add1_dataa <= ( "0000000000000" & Log1p_normal);
	add1 :  prueba1_altfp_log_csa_s0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_add1_dataa,
		datab => almostLog,
		result => wire_add1_result
	  );
	wire_add2_dataa <= ( ER & Log_g(26 DOWNTO 4));
	wire_add2_datab <= ( "000000000000000000000000000000" & round);
	add2 :  prueba1_altfp_log_csa_k0e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_add2_dataa,
		datab => wire_add2_datab,
		result => wire_add2_result
	  );
	exp_biase_sub :  prueba1_altfp_log_csa_0nc
	  PORT MAP ( 
		dataa => exp_data,
		datab => exp_biase,
		result => wire_exp_biase_sub_result
	  );
	wire_sub1_dataa <= (OTHERS => '0');
	sub1 :  prueba1_altfp_log_csa_d4b
	  PORT MAP ( 
		dataa => wire_sub1_dataa,
		datab => Y0(11 DOWNTO 0),
		result => wire_sub1_result
	  );
	wire_sub2_dataa <= (OTHERS => '0');
	sub2 :  prueba1_altfp_log_csa_0nc
	  PORT MAP ( 
		dataa => wire_sub2_dataa,
		datab => E0,
		result => wire_sub2_result
	  );
	wire_sub3_dataa <= ( "0" & lzo);
	wire_sub3_datab <= ( "0" & pfinal_s);
	sub3 :  prueba1_altfp_log_csa_umc
	  PORT MAP ( 
		dataa => wire_sub3_dataa,
		datab => wire_sub3_datab,
		result => wire_sub3_result
	  );
	wire_sub4_datab <= ( "00000000000000" & Z2o2(13 DOWNTO 2));
	sub4 :  prueba1_altfp_log_csa_nlf
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => Zfinal_pipe,
		datab => wire_sub4_datab,
		result => wire_sub4_result
	  );
	wire_sub5_dataa <= ( "0" & "11111" & E0_sub);
	wire_sub5_datab <= ( "000" & lzo_pipe2);
	sub5 :  prueba1_altfp_log_csa_8kf
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => wire_sub5_dataa,
		datab => wire_sub5_datab,
		result => wire_sub5_result
	  );
	wire_sub6_datab <= ( "000" & wire_w_lg_E_normal212w);
	sub6 :  prueba1_altfp_log_csa_0nc
	  PORT MAP ( 
		dataa => E0offset,
		datab => wire_sub6_datab,
		result => wire_sub6_result
	  );
	range_reduction :  prueba1_range_reduction_c2e
	  PORT MAP ( 
		a0_in => man_data(22 DOWNTO 18),
		aclr => aclr,
		almostlog => wire_range_reduction_almostlog,
		clk_en => clk_en,
		clock => clock,
		y0_in => Y0,
		z => wire_range_reduction_z
	  );
	wire_lzc_norm_E_data <= ( Log_normal & "00000000000000001");
	lzc_norm_E :  prueba1_altpriority_encoder_uja
	  PORT MAP ( 
		aclr => aclr,
		clk_en => clk_en,
		clock => clock,
		data => wire_lzc_norm_E_data,
		q => wire_lzc_norm_E_q
	  );
	wire_lzoc_data <= ( wire_w_lg_First_bit96w & "000000001");
	lzoc :  prueba1_altpriority_encoder_q08
	  PORT MAP ( 
		data => wire_lzoc_data,
		q => wire_lzoc_q
	  );
	squarer :  altsquare
	  GENERIC MAP (
		DATA_WIDTH => 13,
		PIPELINE => 1,
		REPRESENTATION => "UNSIGNED",
		RESULT_ALIGNMENT => "MSB",
		RESULT_WIDTH => 14
	  )
	  PORT MAP ( 
		aclr => aclr,
		clock => clock,
		data => squarerIn,
		ena => clk_en,
		result => wire_squarer_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absELog2_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absELog2_pipe_reg0 <= absELog2_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absELog2_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absELog2_pipe_reg1 <= absELog2_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absELog2_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absELog2_pipe_reg2 <= absELog2_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg0 <= absZ0_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg1 <= absZ0_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg2 <= absZ0_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg3 <= absZ0_pipe_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg4 <= absZ0_pipe_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg5 <= absZ0_pipe_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg6 <= absZ0_pipe_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg7 <= absZ0_pipe_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg8 <= absZ0_pipe_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0_pipe_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0_pipe_reg9 <= absZ0_pipe_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0s_pipe1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0s_pipe1_reg0 <= absZ0s_pipe1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0s_pipe1_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0s_pipe1_reg1 <= absZ0s_pipe1_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0s_pipe1_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0s_pipe1_reg2 <= absZ0s_pipe1_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0s_pipe1_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0s_pipe1_reg3 <= absZ0s_pipe1_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN absZ0s_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN absZ0s_reg0 <= absZ0s;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN almostLog_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN almostLog_pipe_reg0 <= almostLog_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN almostLog_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN almostLog_pipe_reg1 <= almostLog_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN almostLog_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN almostLog_pipe_reg2 <= almostLog_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN doRR_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN doRR_reg0(0) <= doRR;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN doRR_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN doRR_reg1 <= doRR_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg0 <= E0_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg1 <= E0_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg2 <= E0_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg3 <= E0_pipe_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg4 <= E0_pipe_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg5 <= E0_pipe_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg6 <= E0_pipe_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg7 <= E0_pipe_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg8 <= E0_pipe_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E0_pipe_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E0_pipe_reg9 <= E0_pipe_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN E_normal_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN E_normal_pipe_reg0 <= E_normal_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_is_ebiase_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_is_ebiase_pipe_reg0(0) <= exp_is_ebiase_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_is_ebiase_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_is_ebiase_pipe_reg1 <= exp_is_ebiase_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_is_ebiase_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_is_ebiase_pipe_reg2 <= exp_is_ebiase_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg0(0) <= input_is_infinity_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg1 <= input_is_infinity_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg10 <= input_is_infinity_pipe_reg9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg11 <= input_is_infinity_pipe_reg10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg12 <= input_is_infinity_pipe_reg11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg13 <= input_is_infinity_pipe_reg12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg14 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg14 <= input_is_infinity_pipe_reg13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg15 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg15 <= input_is_infinity_pipe_reg14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg16 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg16 <= input_is_infinity_pipe_reg15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg17 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg17 <= input_is_infinity_pipe_reg16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg2 <= input_is_infinity_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg3 <= input_is_infinity_pipe_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg4 <= input_is_infinity_pipe_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg5 <= input_is_infinity_pipe_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg6 <= input_is_infinity_pipe_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg7 <= input_is_infinity_pipe_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg8 <= input_is_infinity_pipe_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_infinity_pipe_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_infinity_pipe_reg9 <= input_is_infinity_pipe_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg0(0) <= input_is_nan_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg1 <= input_is_nan_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg10 <= input_is_nan_pipe_reg9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg11 <= input_is_nan_pipe_reg10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg12 <= input_is_nan_pipe_reg11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg13 <= input_is_nan_pipe_reg12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg14 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg14 <= input_is_nan_pipe_reg13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg15 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg15 <= input_is_nan_pipe_reg14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg16 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg16 <= input_is_nan_pipe_reg15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg17 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg17 <= input_is_nan_pipe_reg16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg2 <= input_is_nan_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg3 <= input_is_nan_pipe_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg4 <= input_is_nan_pipe_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg5 <= input_is_nan_pipe_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg6 <= input_is_nan_pipe_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg7 <= input_is_nan_pipe_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg8 <= input_is_nan_pipe_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_nan_pipe_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_nan_pipe_reg9 <= input_is_nan_pipe_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg0(0) <= input_is_one_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg1 <= input_is_one_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg10 <= input_is_one_pipe_reg9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg11 <= input_is_one_pipe_reg10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg12 <= input_is_one_pipe_reg11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg13 <= input_is_one_pipe_reg12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg14 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg14 <= input_is_one_pipe_reg13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg15 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg15 <= input_is_one_pipe_reg14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg16 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg16 <= input_is_one_pipe_reg15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg17 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg17 <= input_is_one_pipe_reg16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg2 <= input_is_one_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg3 <= input_is_one_pipe_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg4 <= input_is_one_pipe_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg5 <= input_is_one_pipe_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg6 <= input_is_one_pipe_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg7 <= input_is_one_pipe_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg8 <= input_is_one_pipe_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_one_pipe_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_one_pipe_reg9 <= input_is_one_pipe_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg0(0) <= input_is_zero_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg1 <= input_is_zero_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg10 <= input_is_zero_pipe_reg9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg11 <= input_is_zero_pipe_reg10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg12 <= input_is_zero_pipe_reg11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg13 <= input_is_zero_pipe_reg12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg14 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg14 <= input_is_zero_pipe_reg13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg15 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg15 <= input_is_zero_pipe_reg14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg16 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg16 <= input_is_zero_pipe_reg15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg17 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg17 <= input_is_zero_pipe_reg16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg2 <= input_is_zero_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg3 <= input_is_zero_pipe_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg4 <= input_is_zero_pipe_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg5 <= input_is_zero_pipe_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg6 <= input_is_zero_pipe_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg7 <= input_is_zero_pipe_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg8 <= input_is_zero_pipe_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_is_zero_pipe_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_is_zero_pipe_reg9 <= input_is_zero_pipe_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Log_normal_normd_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Log_normal_normd_pipe_reg0 <= Log_normal_normd_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Log_normal_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Log_normal_reg0 <= Log_normal;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Log_small_normd_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Log_small_normd_pipe_reg0 <= Log_small_normd_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Log_small_normd_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Log_small_normd_pipe_reg1 <= Log_small_normd_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Lshiftval_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Lshiftval_reg0 <= Lshiftval;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Lshiftval_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Lshiftval_reg1 <= Lshiftval_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Lshiftval_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Lshiftval_reg2 <= Lshiftval_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Lshiftval_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Lshiftval_reg3 <= Lshiftval_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg0 <= lzo_pipe1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg1 <= lzo_pipe1_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg2 <= lzo_pipe1_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg3 <= lzo_pipe1_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg4 <= lzo_pipe1_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg5 <= lzo_pipe1_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg6 <= lzo_pipe1_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg7 <= lzo_pipe1_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg8 <= lzo_pipe1_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_pipe1_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_pipe1_reg9 <= lzo_pipe1_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg0 <= lzo;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg1 <= lzo_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg2 <= lzo_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg3 <= lzo_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg4 <= lzo_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg5 <= lzo_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg6 <= lzo_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN lzo_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN lzo_reg7 <= lzo_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_data_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_data_reg0(0) <= sign_data;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_data_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_data_reg1 <= sign_data_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_data_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_data_reg2 <= sign_data_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg0(0) <= small_flag_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg1 <= small_flag_pipe_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg2 <= small_flag_pipe_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg3 <= small_flag_pipe_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg4 <= small_flag_pipe_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg5 <= small_flag_pipe_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg6 <= small_flag_pipe_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg7 <= small_flag_pipe_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg8 <= small_flag_pipe_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN small_flag_pipe_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN small_flag_pipe_reg9 <= small_flag_pipe_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg0(0) <= sR_pipe1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg1 <= sR_pipe1_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg2 <= sR_pipe1_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg3 <= sR_pipe1_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg4 <= sR_pipe1_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg5 <= sR_pipe1_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg6 <= sR_pipe1_reg5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg7 <= sR_pipe1_reg6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg8 <= sR_pipe1_reg7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe1_reg9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe1_reg9 <= sR_pipe1_reg8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe2_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe2_reg0(0) <= sR_pipe2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe2_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe2_reg1 <= sR_pipe2_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe2_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe2_reg2 <= sR_pipe2_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe2_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe2_reg3 <= sR_pipe2_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe2_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe2_reg4 <= sR_pipe2_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe2_reg5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe2_reg5 <= sR_pipe2_reg4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe3_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe3_reg0(0) <= sR_pipe3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe3_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe3_reg1 <= sR_pipe3_reg0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe3_reg2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe3_reg2 <= sR_pipe3_reg1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe3_reg3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe3_reg3 <= sR_pipe3_reg2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sR_pipe3_reg4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sR_pipe3_reg4 <= sR_pipe3_reg3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Z2o2_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Z2o2_pipe_reg0 <= Z2o2_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Z2o2_small_s_pipe_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Z2o2_small_s_pipe_reg0 <= Z2o2_small_s_pipe;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Zfinal_reg0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Zfinal_reg0 <= Zfinal;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Zfinal_reg1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN Zfinal_reg1 <= Zfinal_reg0;
			END IF;
		END IF;
	END PROCESS;
	addsub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_PIPELINE => 2,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 29
	  )
	  PORT MAP ( 
		add_sub => sR_pipe3,
		clock => clock,
		dataa => Z_small,
		datab => Z2o2_small,
		result => wire_addsub1_result
	  );
	wire_addsub2_add_sub <= wire_w_lg_sR_pipe3179w(0);
	addsub2 :  lpm_add_sub
	  GENERIC MAP (
		LPM_PIPELINE => 2,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 47
	  )
	  PORT MAP ( 
		add_sub => wire_addsub2_add_sub,
		clock => clock,
		dataa => absELog2_pad,
		datab => LogF_normal_pad,
		result => wire_addsub2_result
	  );
	mult1 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 8,
		LPM_WIDTHB => 27,
		LPM_WIDTHP => 35
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => absE,
		datab => Log2,
		result => wire_mult1_result
	  );
	wire_mux_result0a_dataout <= ( wire_w_lg_w_lg_input_is_one247w248w & wire_w_lg_w_lg_input_is_one247w248w & wire_w_lg_w_lg_input_is_one247w248w & wire_w_lg_w_lg_input_is_one247w248w & wire_w_lg_w_lg_input_is_one247w248w & wire_w_lg_w_lg_input_is_one247w248w & wire_w_lg_w_lg_input_is_one247w248w & wire_w_lg_w_lg_input_is_one247w248w & input_is_nan & "0000000000000000000000") WHEN wire_w_lg_w_lg_w_lg_input_is_zero244w245w246w(0) = '1'  ELSE EFR;

 END RTL; --prueba1_altfp_log_8ka
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY prueba1 IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END prueba1;


ARCHITECTURE RTL OF prueba1 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT prueba1_altfp_log_8ka
	PORT (
			clock	: IN STD_LOGIC ;
			data	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	prueba1_altfp_log_8ka_component : prueba1_altfp_log_8ka
	PORT MAP (
		clock => clock,
		data => data,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altfp_log"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "21"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: USED_PORT: data 0 0 32 0 INPUT NODEFVAL "data[31..0]"
-- Retrieval info: CONNECT: @data 0 0 32 0 data 0 0 32 0
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL prueba1.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL prueba1.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL prueba1.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL prueba1_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL prueba1.inc FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL prueba1.cmp TRUE TRUE
-- Retrieval info: LIB_FILE: lpm
